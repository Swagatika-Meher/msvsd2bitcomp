MACRO 1BITADC
  ORIGIN 0 0 ;
  FOREIGN 1BITADC 0 0 ;
  SIZE 11.18 BY 15.12 ;
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 6.58 2.32 6.86 ;
      LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
      LAYER M2 ;
        RECT 1.56 6.58 1.88 6.86 ;
      LAYER M3 ;
        RECT 1.58 6.72 1.86 7.98 ;
      LAYER M2 ;
        RECT 1.56 7.84 1.88 8.12 ;
    END
  END OUT
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 1.15 0.68 1.43 6.46 ;
      LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
      LAYER M3 ;
        RECT 1.15 3.595 1.43 3.965 ;
      LAYER M2 ;
        RECT 1.29 3.64 4.3 3.92 ;
      LAYER M3 ;
        RECT 4.16 3.595 4.44 3.965 ;
      LAYER M2 ;
        RECT 6.28 0.7 7.48 0.98 ;
      LAYER M3 ;
        RECT 4.16 1.075 4.44 1.445 ;
      LAYER M2 ;
        RECT 4.3 1.12 6.02 1.4 ;
      LAYER M1 ;
        RECT 5.895 0.84 6.145 1.26 ;
      LAYER M2 ;
        RECT 6.02 0.7 6.45 0.98 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 0.72 8.24 1 14.44 ;
      LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
      LAYER M3 ;
        RECT 6.31 8.66 6.59 14.44 ;
      LAYER M3 ;
        RECT 0.72 11.155 1 11.525 ;
      LAYER M2 ;
        RECT 0.86 11.2 4.3 11.48 ;
      LAYER M3 ;
        RECT 4.16 11.155 4.44 11.525 ;
      LAYER M2 ;
        RECT 4.3 11.2 6.45 11.48 ;
      LAYER M3 ;
        RECT 6.31 11.155 6.59 11.525 ;
    END
  END VDD
  PIN INP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.86 4.06 10.06 4.34 ;
    END
  END INP
  PIN INN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
    END
  END INN
  OBS 
  LAYER M3 ;
        RECT 2.01 2.78 2.29 7.3 ;
  LAYER M2 ;
        RECT 4.56 2.8 5.76 3.08 ;
  LAYER M3 ;
        RECT 2.01 3.175 2.29 3.545 ;
  LAYER M2 ;
        RECT 2.15 3.22 3.87 3.5 ;
  LAYER M1 ;
        RECT 3.745 2.94 3.995 3.36 ;
  LAYER M2 ;
        RECT 3.87 2.8 4.73 3.08 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 12.34 ;
  LAYER M3 ;
        RECT 2.01 7.14 2.29 7.56 ;
  LAYER M2 ;
        RECT 2.15 7.42 3.87 7.7 ;
  LAYER M3 ;
        RECT 3.73 7.56 4.01 7.98 ;
  LAYER M2 ;
        RECT 1.99 7.42 2.31 7.7 ;
  LAYER M3 ;
        RECT 2.01 7.4 2.29 7.72 ;
  LAYER M2 ;
        RECT 3.71 7.42 4.03 7.7 ;
  LAYER M3 ;
        RECT 3.73 7.4 4.01 7.72 ;
  LAYER M2 ;
        RECT 1.99 7.42 2.31 7.7 ;
  LAYER M3 ;
        RECT 2.01 7.4 2.29 7.72 ;
  LAYER M2 ;
        RECT 3.71 7.42 4.03 7.7 ;
  LAYER M3 ;
        RECT 3.73 7.4 4.01 7.72 ;
  LAYER M2 ;
        RECT 4.56 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 6.71 6.58 7.91 6.86 ;
  LAYER M3 ;
        RECT 10.18 1.94 10.46 8.14 ;
  LAYER M2 ;
        RECT 5.43 7 5.75 7.28 ;
  LAYER M1 ;
        RECT 5.465 6.3 5.715 7.14 ;
  LAYER M2 ;
        RECT 5.59 6.16 6.88 6.44 ;
  LAYER M3 ;
        RECT 6.74 6.3 7.02 6.72 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M2 ;
        RECT 7.74 6.58 10.32 6.86 ;
  LAYER M3 ;
        RECT 10.18 6.535 10.46 6.905 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 5.465 7.055 5.715 7.225 ;
  LAYER M2 ;
        RECT 5.42 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 6.72 6.16 7.04 6.44 ;
  LAYER M3 ;
        RECT 6.74 6.14 7.02 6.46 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 5.465 7.055 5.715 7.225 ;
  LAYER M2 ;
        RECT 5.42 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 6.72 6.16 7.04 6.44 ;
  LAYER M3 ;
        RECT 6.74 6.14 7.02 6.46 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 5.465 7.055 5.715 7.225 ;
  LAYER M2 ;
        RECT 5.42 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 6.72 6.16 7.04 6.44 ;
  LAYER M3 ;
        RECT 6.74 6.14 7.02 6.46 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M2 ;
        RECT 10.16 6.58 10.48 6.86 ;
  LAYER M3 ;
        RECT 10.18 6.56 10.46 6.88 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 5.465 7.055 5.715 7.225 ;
  LAYER M2 ;
        RECT 5.42 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 6.72 6.16 7.04 6.44 ;
  LAYER M3 ;
        RECT 6.74 6.14 7.02 6.46 ;
  LAYER M2 ;
        RECT 6.72 6.58 7.04 6.86 ;
  LAYER M3 ;
        RECT 6.74 6.56 7.02 6.88 ;
  LAYER M2 ;
        RECT 10.16 6.58 10.48 6.86 ;
  LAYER M3 ;
        RECT 10.18 6.56 10.46 6.88 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 12.34 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 7.14 7.45 7.98 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 6.98 7.45 7.3 ;
  LAYER M2 ;
        RECT 7.15 7 7.47 7.28 ;
  LAYER M3 ;
        RECT 7.17 6.98 7.45 7.3 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 6.28 8.26 7.48 8.54 ;
  LAYER M2 ;
        RECT 8.86 8.26 10.06 8.54 ;
  LAYER M2 ;
        RECT 1.99 12.04 2.31 12.32 ;
  LAYER M1 ;
        RECT 2.025 9.24 2.275 12.18 ;
  LAYER M2 ;
        RECT 2.15 9.1 6.02 9.38 ;
  LAYER M3 ;
        RECT 5.88 8.4 6.16 9.24 ;
  LAYER M2 ;
        RECT 6.02 8.26 6.45 8.54 ;
  LAYER M2 ;
        RECT 7.31 8.26 9.03 8.54 ;
  LAYER M1 ;
        RECT 2.025 9.155 2.275 9.325 ;
  LAYER M2 ;
        RECT 1.98 9.1 2.32 9.38 ;
  LAYER M1 ;
        RECT 2.025 12.095 2.275 12.265 ;
  LAYER M2 ;
        RECT 1.98 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 5.86 8.26 6.18 8.54 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 8.56 ;
  LAYER M2 ;
        RECT 5.86 9.1 6.18 9.38 ;
  LAYER M3 ;
        RECT 5.88 9.08 6.16 9.4 ;
  LAYER M1 ;
        RECT 2.025 9.155 2.275 9.325 ;
  LAYER M2 ;
        RECT 1.98 9.1 2.32 9.38 ;
  LAYER M1 ;
        RECT 2.025 12.095 2.275 12.265 ;
  LAYER M2 ;
        RECT 1.98 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 5.86 8.26 6.18 8.54 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 8.56 ;
  LAYER M2 ;
        RECT 5.86 9.1 6.18 9.38 ;
  LAYER M3 ;
        RECT 5.88 9.08 6.16 9.4 ;
  LAYER M1 ;
        RECT 2.025 9.155 2.275 9.325 ;
  LAYER M2 ;
        RECT 1.98 9.1 2.32 9.38 ;
  LAYER M1 ;
        RECT 2.025 12.095 2.275 12.265 ;
  LAYER M2 ;
        RECT 1.98 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 5.86 8.26 6.18 8.54 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 8.56 ;
  LAYER M2 ;
        RECT 5.86 9.1 6.18 9.38 ;
  LAYER M3 ;
        RECT 5.88 9.08 6.16 9.4 ;
  LAYER M1 ;
        RECT 2.025 9.155 2.275 9.325 ;
  LAYER M2 ;
        RECT 1.98 9.1 2.32 9.38 ;
  LAYER M1 ;
        RECT 2.025 12.095 2.275 12.265 ;
  LAYER M2 ;
        RECT 1.98 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 5.86 8.26 6.18 8.54 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 8.56 ;
  LAYER M2 ;
        RECT 5.86 9.1 6.18 9.38 ;
  LAYER M3 ;
        RECT 5.88 9.08 6.16 9.4 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
  LAYER M2 ;
        RECT 1.98 7 3.18 7.28 ;
  LAYER M2 ;
        RECT 0.69 6.16 2.75 6.44 ;
  LAYER M2 ;
        RECT 1.12 0.7 2.32 0.98 ;
  LAYER M3 ;
        RECT 2.01 2.78 2.29 7.3 ;
  LAYER M2 ;
        RECT 1.12 6.58 2.32 6.86 ;
  LAYER M3 ;
        RECT 1.15 0.68 1.43 6.46 ;
  LAYER M1 ;
        RECT 4.605 3.695 4.855 7.225 ;
  LAYER M1 ;
        RECT 4.605 2.435 4.855 3.445 ;
  LAYER M1 ;
        RECT 4.605 0.335 4.855 1.345 ;
  LAYER M1 ;
        RECT 5.035 3.695 5.285 7.225 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M2 ;
        RECT 4.13 6.58 5.33 6.86 ;
  LAYER M2 ;
        RECT 4.13 0.7 5.33 0.98 ;
  LAYER M2 ;
        RECT 4.56 7 5.76 7.28 ;
  LAYER M2 ;
        RECT 4.56 2.8 5.76 3.08 ;
  LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 11.425 ;
  LAYER M1 ;
        RECT 7.185 11.675 7.435 12.685 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 14.785 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M2 ;
        RECT 7.14 7.84 8.34 8.12 ;
  LAYER M2 ;
        RECT 5.85 8.68 7.91 8.96 ;
  LAYER M2 ;
        RECT 6.28 14.14 7.48 14.42 ;
  LAYER M3 ;
        RECT 7.17 7.82 7.45 12.34 ;
  LAYER M2 ;
        RECT 6.28 8.26 7.48 8.54 ;
  LAYER M3 ;
        RECT 6.31 8.66 6.59 14.44 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 2.84 12.04 4.04 12.32 ;
  LAYER M2 ;
        RECT 2.84 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 12.34 ;
  LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
  LAYER M1 ;
        RECT 9.765 4.955 10.015 8.485 ;
  LAYER M1 ;
        RECT 9.765 3.695 10.015 4.705 ;
  LAYER M1 ;
        RECT 9.765 1.595 10.015 2.605 ;
  LAYER M1 ;
        RECT 9.335 4.955 9.585 8.485 ;
  LAYER M1 ;
        RECT 10.195 4.955 10.445 8.485 ;
  LAYER M2 ;
        RECT 9.29 7.84 10.49 8.12 ;
  LAYER M2 ;
        RECT 9.29 1.96 10.49 2.24 ;
  LAYER M2 ;
        RECT 8.86 8.26 10.06 8.54 ;
  LAYER M2 ;
        RECT 8.86 4.06 10.06 4.34 ;
  LAYER M3 ;
        RECT 10.18 1.94 10.46 8.14 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M3 ;
        RECT 0.72 8.24 1 14.44 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M2 ;
        RECT 6.28 0.7 7.48 0.98 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 6.71 6.58 7.91 6.86 ;
  END 
END 1BITADC
