** sch_path: /home/swagatika/Desktop/Circuits/1_bit_ADC_sym.sch
.subckt 1_bit_ADC_sym Vdd INN INP Gnd OUT
*.PININFO Vdd:B INN:B INP:B Gnd:B OUT:O
XM2 net1 net3 Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 net3 INN net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net1 INP net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM1 net3 net3 Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 OUT net1 Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 OUT net4 Gnd Gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM7 net2 net4 Gnd Gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 net4 net4 Gnd Gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM9 net4 net4 Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
.ends
.end
