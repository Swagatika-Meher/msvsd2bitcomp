* SPICE3 file created from INVERTER_0.ext - technology: sky130A

X0 OUT IN GND GND sky130_fd_pr__nfet_01v8 ad=2.94e+11p pd=2.66e+06u as=5.565e+11p ps=5.26e+06u w=1.05e+06u l=150000u
X1 GND IN OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X2 OUT IN INV_33483112_0_0_1676996573_0/PMOS_S_3683112_X1_Y1_1676996573_1676996573_0/w_0_0# INV_33483112_0_0_1676996573_0/PMOS_S_3683112_X1_Y1_1676996573_1676996573_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=2.94e+11p pd=2.66e+06u as=5.565e+11p ps=5.26e+06u w=1.05e+06u l=150000u
X3 INV_33483112_0_0_1676996573_0/PMOS_S_3683112_X1_Y1_1676996573_1676996573_0/w_0_0# IN OUT INV_33483112_0_0_1676996573_0/PMOS_S_3683112_X1_Y1_1676996573_1676996573_0/w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
C0 IN INV_33483112_0_0_1676996573_0/PMOS_S_3683112_X1_Y1_1676996573_1676996573_0/w_0_0# 1.10fF
C1 OUT INV_33483112_0_0_1676996573_0/PMOS_S_3683112_X1_Y1_1676996573_1676996573_0/w_0_0# 0.79fF
C2 IN OUT 0.31fF
C3 OUT GND 0.69fF **FLOATING
C4 IN GND 1.45fF **FLOATING
C5 INV_33483112_0_0_1676996573_0/PMOS_S_3683112_X1_Y1_1676996573_1676996573_0/w_0_0# GND 3.02fF **FLOATING
