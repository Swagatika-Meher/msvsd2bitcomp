magic
tech sky130A
magscale 1 2
timestamp 1676651141
<< metal1 >>
rect -7252 1082 -6838 1084
rect -7296 1076 -6754 1082
rect -3404 1076 -3204 1224
rect -7296 1072 -1256 1076
rect -7296 974 1742 1072
rect -7296 972 -6754 974
rect -7296 970 -6894 972
rect -7296 112 -7212 970
rect -6854 190 -6792 248
rect -5562 186 -5498 244
rect -4176 196 -4116 252
rect -2456 188 -2394 248
rect -692 212 -634 268
rect 908 220 966 282
rect 1496 154 1736 974
rect -638 148 894 152
rect -2114 130 -1980 132
rect -6022 126 -5930 130
rect -7296 -26 -6856 112
rect -6798 -26 -5562 126
rect -5500 116 -5056 118
rect -4868 116 -4604 118
rect -4502 116 -4176 118
rect -5500 102 -4176 116
rect -5500 16 -5022 102
rect -4902 16 -4176 102
rect -5500 -8 -4176 16
rect -5500 -14 -5056 -8
rect -4868 -14 -4176 -8
rect -4122 110 -2456 130
rect -4122 2 -3302 110
rect -3186 2 -2456 110
rect -4122 -24 -2456 2
rect -2390 116 -694 130
rect -2390 20 -1588 116
rect -1368 20 -694 116
rect -638 24 908 148
rect -638 22 894 24
rect -2390 2 -694 20
rect 964 10 1736 154
rect 1496 2 1736 10
rect -2390 -4 -1622 2
rect -1334 -4 -694 2
rect -7296 -36 -7212 -26
rect -4122 -28 -3328 -24
rect -3162 -28 -2456 -24
rect -6858 -522 -6788 -88
rect -5562 -522 -5502 -90
rect -4174 -506 -4118 -82
rect -2452 -482 -2402 -88
rect -688 -478 -632 -64
rect -6926 -722 -6726 -522
rect -5640 -722 -5440 -522
rect -4244 -706 -4044 -506
rect -2530 -682 -2330 -482
rect -756 -678 -556 -478
rect 908 -482 964 -58
rect -6868 -1116 -6798 -722
rect -7200 -1252 -6796 -1116
rect -7196 -2080 -7126 -1252
rect -5560 -2064 -5504 -722
rect -4178 -2060 -4124 -706
rect -3302 -1092 -3204 -1082
rect -3302 -1200 -3296 -1092
rect -3210 -1200 -3204 -1092
rect -3302 -1440 -3204 -1200
rect -3336 -1640 -3136 -1440
rect -2460 -2040 -2410 -682
rect -696 -2034 -646 -678
rect 852 -682 1052 -482
rect 898 -2020 954 -682
rect -2410 -2092 -1936 -2088
rect -4600 -2126 -4186 -2106
rect -7622 -2140 -7568 -2136
rect -7132 -2140 -6470 -2138
rect -6134 -2140 -5566 -2138
rect -7622 -2150 -7190 -2140
rect -7622 -2280 -7606 -2150
rect -7542 -2280 -7190 -2150
rect -7132 -2156 -5566 -2140
rect -7132 -2236 -6440 -2156
rect -6184 -2236 -5566 -2156
rect -7132 -2264 -5566 -2236
rect -7132 -2266 -6470 -2264
rect -7132 -2270 -6826 -2266
rect -6706 -2270 -6470 -2266
rect -6134 -2270 -5566 -2264
rect -5504 -2142 -5018 -2128
rect -5504 -2262 -5084 -2142
rect -5032 -2262 -5018 -2142
rect -5504 -2278 -5018 -2262
rect -4600 -2260 -4584 -2126
rect -4502 -2260 -4186 -2126
rect -4122 -2246 -2462 -2112
rect -2410 -2242 -1882 -2092
rect -4122 -2248 -3804 -2246
rect -3660 -2248 -2462 -2246
rect -4600 -2278 -4186 -2260
rect -5504 -2280 -5022 -2278
rect -7622 -2294 -7190 -2280
rect -7622 -2296 -7568 -2294
rect -7190 -2346 -7130 -2344
rect -7192 -2400 -7130 -2346
rect -5566 -2386 -5504 -2330
rect -4186 -2380 -4122 -2322
rect -2466 -2356 -2404 -2300
rect -7190 -2402 -7130 -2400
rect -2012 -3068 -1882 -2242
rect -1136 -2248 -706 -2084
rect -646 -2104 894 -2084
rect -646 -2200 -14 -2104
rect 162 -2200 894 -2104
rect -646 -2226 894 -2200
rect 952 -2222 1352 -2084
rect -646 -2228 -40 -2226
rect 192 -2228 894 -2226
rect -1136 -3068 -1024 -2248
rect 894 -2280 954 -2278
rect -704 -2352 -640 -2300
rect 894 -2332 956 -2280
rect -712 -3068 -626 -3066
rect 878 -3068 984 -3064
rect 1288 -3068 1352 -2222
rect -2016 -3198 1352 -3068
rect -2016 -3208 1348 -3198
rect -2016 -3212 978 -3208
rect -722 -3304 -632 -3212
rect -766 -3504 -566 -3304
<< via1 >>
rect -5022 16 -4902 102
rect -3302 2 -3186 110
rect -1588 20 -1368 116
rect -3296 -1200 -3210 -1092
rect -7606 -2280 -7542 -2150
rect -6440 -2236 -6184 -2156
rect -5084 -2262 -5032 -2142
rect -4584 -2260 -4502 -2126
rect -14 -2200 162 -2104
<< metal2 >>
rect -5034 764 -1508 768
rect -5034 722 -1348 764
rect -5036 686 -1348 722
rect -5036 272 -4884 686
rect -5036 102 -4882 272
rect -1612 252 -1348 686
rect -5036 16 -5022 102
rect -4902 16 -4882 102
rect -5036 -8 -4882 16
rect -3328 110 -3162 146
rect -3328 2 -3302 110
rect -3186 2 -3162 110
rect -3328 -60 -3162 2
rect -1614 116 -1344 252
rect -1614 20 -1588 116
rect -1368 20 -1344 116
rect -1614 -4 -1344 20
rect -5930 -1078 -5816 -1076
rect -3302 -1078 -3196 -60
rect -5930 -1092 -3196 -1078
rect -5930 -1200 -3296 -1092
rect -3210 -1200 -3196 -1092
rect -5930 -1210 -3198 -1200
rect -7594 -1442 -7410 -1440
rect -7596 -1446 -7410 -1442
rect -5930 -1446 -5816 -1210
rect -7596 -1540 -5816 -1446
rect -7596 -2136 -7530 -1540
rect -7484 -1542 -5816 -1540
rect -5930 -1550 -5816 -1542
rect -5096 -2126 -5014 -1210
rect -7622 -2140 -7530 -2136
rect -7622 -2150 -7528 -2140
rect -7622 -2280 -7606 -2150
rect -7542 -2280 -7528 -2150
rect -7622 -2296 -7528 -2280
rect -6472 -2156 -6150 -2140
rect -6472 -2236 -6440 -2156
rect -6184 -2236 -6150 -2156
rect -6472 -2304 -6150 -2236
rect -5092 -2142 -5014 -2126
rect -5092 -2262 -5084 -2142
rect -5032 -2262 -5014 -2142
rect -5092 -2276 -5014 -2262
rect -4606 -2122 -4484 -1210
rect -40 -2104 190 -2080
rect -4606 -2126 -4482 -2122
rect -4606 -2260 -4584 -2126
rect -4502 -2260 -4482 -2126
rect -4606 -2276 -4482 -2260
rect -40 -2200 -14 -2104
rect 162 -2200 190 -2104
rect -5092 -2284 -5018 -2276
rect -6472 -2340 -6148 -2304
rect -6464 -3528 -6148 -2340
rect -6464 -3574 -6152 -3528
rect -40 -3536 190 -2200
rect -6462 -3600 -6152 -3574
rect -42 -3600 196 -3536
rect -6462 -3734 196 -3600
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1676639765
transform 1 0 -6823 0 1 49
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM2
timestamp 1676639765
transform 1 0 937 0 1 81
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3
timestamp 1676639765
transform 1 0 -5529 0 1 47
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM4
timestamp 1676639765
transform 1 0 -661 0 1 73
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM5
timestamp 1676639765
transform 1 0 -4145 0 1 55
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM6
timestamp 1676639765
transform 1 0 -2423 0 1 51
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM7
timestamp 1676639765
transform 1 0 -7161 0 1 -2216
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM8
timestamp 1676639765
transform 1 0 -5535 0 1 -2202
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM9
timestamp 1676639765
transform 1 0 -4153 0 1 -2194
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM10
timestamp 1676639765
transform 1 0 925 0 1 -2150
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM11
timestamp 1676639765
transform 1 0 -673 0 1 -2168
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM12
timestamp 1676639765
transform 1 0 -2435 0 1 -2172
box -211 -310 211 310
<< labels >>
flabel metal1 -3404 1024 -3204 1224 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -5640 -722 -5440 -522 0 FreeSans 256 0 0 0 C
port 4 nsew
flabel metal1 -4244 -706 -4044 -506 0 FreeSans 256 0 0 0 E
port 6 nsew
flabel metal1 -2530 -682 -2330 -482 0 FreeSans 256 0 0 0 F
port 5 nsew
flabel metal1 -756 -678 -556 -478 0 FreeSans 256 0 0 0 D
port 3 nsew
flabel metal1 852 -682 1052 -482 0 FreeSans 256 0 0 0 B
port 2 nsew
flabel metal1 -6926 -722 -6726 -522 0 FreeSans 256 0 0 0 A
port 1 nsew
flabel metal1 -766 -3504 -566 -3304 0 FreeSans 256 0 0 0 Gnd
port 8 nsew
flabel metal1 -3336 -1640 -3136 -1440 0 FreeSans 256 0 0 0 Fn
port 7 nsew
<< end >>
