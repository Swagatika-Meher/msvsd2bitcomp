magic
tech sky130A
magscale 1 2
timestamp 1677569328
<< nwell >>
rect 0 0 516 1512
<< pmos >>
rect 200 462 230 672
rect 286 462 316 672
<< pdiff >>
rect 147 648 200 672
rect 147 614 155 648
rect 189 614 200 648
rect 147 580 200 614
rect 147 546 155 580
rect 189 546 200 580
rect 147 512 200 546
rect 147 478 155 512
rect 189 478 200 512
rect 147 462 200 478
rect 230 648 286 672
rect 230 614 241 648
rect 275 614 286 648
rect 230 580 286 614
rect 230 546 241 580
rect 275 546 286 580
rect 230 512 286 546
rect 230 478 241 512
rect 275 478 286 512
rect 230 462 286 478
rect 316 648 369 672
rect 316 614 327 648
rect 361 614 369 648
rect 316 580 369 614
rect 316 546 327 580
rect 361 546 369 580
rect 316 512 369 546
rect 316 478 327 512
rect 361 478 369 512
rect 316 462 369 478
<< pdiffc >>
rect 155 614 189 648
rect 155 546 189 580
rect 155 478 189 512
rect 241 614 275 648
rect 241 546 275 580
rect 241 478 275 512
rect 327 614 361 648
rect 327 546 361 580
rect 327 478 361 512
<< nsubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
<< nsubdiffcont >>
rect 241 1327 275 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 672 230 897
rect 286 672 316 897
rect 200 252 230 462
rect 286 252 316 462
<< polycont >>
rect 241 907 275 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 147 648 197 773
rect 147 614 155 648
rect 189 614 197 648
rect 147 580 197 614
rect 147 546 155 580
rect 189 546 197 580
rect 147 512 197 546
rect 147 478 155 512
rect 189 478 197 512
rect 147 185 197 478
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 648 283 773
rect 233 614 241 648
rect 275 614 283 648
rect 233 580 283 614
rect 233 546 241 580
rect 275 546 283 580
rect 233 512 283 546
rect 233 478 241 512
rect 275 478 283 512
rect 233 101 283 478
rect 233 67 241 101
rect 275 67 283 101
rect 319 648 369 773
rect 319 614 327 648
rect 361 614 369 648
rect 319 580 369 614
rect 319 546 327 580
rect 361 546 369 580
rect 319 512 369 546
rect 319 478 327 512
rect 361 478 369 512
rect 319 185 369 478
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
<< viali >>
rect 241 1327 275 1361
rect 241 907 275 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
<< metal1 >>
rect 138 1370 378 1372
rect 138 1361 318 1370
rect 138 1327 241 1361
rect 275 1327 318 1361
rect 138 1318 318 1327
rect 370 1318 378 1370
rect 138 1316 378 1318
rect 52 941 292 952
rect 52 907 241 941
rect 275 907 292 941
rect 52 896 292 907
rect 138 194 378 196
rect 138 185 318 194
rect 138 151 155 185
rect 189 151 318 185
rect 138 142 318 151
rect 370 142 378 194
rect 138 140 378 142
rect 52 101 292 112
rect 52 67 241 101
rect 275 67 292 101
rect 52 56 292 67
<< via1 >>
rect 318 1318 370 1370
rect 318 185 370 194
rect 318 151 327 185
rect 327 151 361 185
rect 361 151 370 185
rect 318 142 370 151
<< metal2 >>
rect 316 1370 372 1376
rect 316 1318 318 1370
rect 370 1318 372 1370
rect 316 194 372 1318
rect 316 142 318 194
rect 370 142 372 194
rect 316 136 372 142
<< end >>
