MACRO RINGOSCILLATOR
  ORIGIN 0 0 ;
  FOREIGN RINGOSCILLATOR 0 0 ;
  SIZE 10.32 BY 30.24 ;
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 2.87 8.24 3.15 14.44 ;
      LAYER M3 ;
        RECT 7.17 8.24 7.45 14.44 ;
      LAYER M3 ;
        RECT 2.87 11.155 3.15 11.525 ;
      LAYER M2 ;
        RECT 3.01 11.2 7.31 11.48 ;
      LAYER M3 ;
        RECT 7.17 11.155 7.45 11.525 ;
      LAYER M3 ;
        RECT 4.59 23.36 4.87 29.56 ;
      LAYER M3 ;
        RECT 2.87 14.28 3.15 22.68 ;
      LAYER M2 ;
        RECT 3.01 22.54 4.73 22.82 ;
      LAYER M3 ;
        RECT 4.59 22.68 4.87 23.52 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 2.87 0.68 3.15 6.88 ;
      LAYER M3 ;
        RECT 7.17 0.68 7.45 6.88 ;
      LAYER M3 ;
        RECT 2.87 3.595 3.15 3.965 ;
      LAYER M2 ;
        RECT 3.01 3.64 7.31 3.92 ;
      LAYER M3 ;
        RECT 7.17 3.595 7.45 3.965 ;
      LAYER M3 ;
        RECT 4.59 15.8 4.87 22 ;
      LAYER M3 ;
        RECT 7.17 6.72 7.45 7.56 ;
      LAYER M2 ;
        RECT 6.88 7.42 7.31 7.7 ;
      LAYER M3 ;
        RECT 6.74 7.56 7.02 14.7 ;
      LAYER M2 ;
        RECT 4.73 14.56 6.88 14.84 ;
      LAYER M3 ;
        RECT 4.59 14.7 4.87 15.96 ;
    END
  END VDD
  PIN OUT
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 1.12 2.8 4.04 3.08 ;
      LAYER M2 ;
        RECT 1.12 12.04 4.04 12.32 ;
      LAYER M2 ;
        RECT 2.42 2.8 2.74 3.08 ;
      LAYER M3 ;
        RECT 2.44 2.94 2.72 12.18 ;
      LAYER M2 ;
        RECT 2.42 12.04 2.74 12.32 ;
      LAYER M2 ;
        RECT 3.7 22.12 6.62 22.4 ;
      LAYER M2 ;
        RECT 3.7 22.96 6.62 23.24 ;
      LAYER M2 ;
        RECT 5 22.12 5.32 22.4 ;
      LAYER M3 ;
        RECT 5.02 22.26 5.3 23.1 ;
      LAYER M2 ;
        RECT 5 22.96 5.32 23.24 ;
      LAYER M2 ;
        RECT 3.71 12.04 4.03 12.32 ;
      LAYER M3 ;
        RECT 3.73 12.18 4.01 22.26 ;
      LAYER M2 ;
        RECT 3.71 22.12 4.03 22.4 ;
    END
  END OUT
  OBS 
  LAYER M2 ;
        RECT 6.28 7 9.2 7.28 ;
  LAYER M2 ;
        RECT 6.28 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 7.58 7 7.9 7.28 ;
  LAYER M3 ;
        RECT 7.6 7.14 7.88 7.98 ;
  LAYER M2 ;
        RECT 7.58 7.84 7.9 8.12 ;
  LAYER M2 ;
        RECT 3.7 17.92 6.62 18.2 ;
  LAYER M2 ;
        RECT 3.7 27.16 6.62 27.44 ;
  LAYER M2 ;
        RECT 5.43 17.92 5.75 18.2 ;
  LAYER M3 ;
        RECT 5.45 18.06 5.73 27.3 ;
  LAYER M2 ;
        RECT 5.43 27.16 5.75 27.44 ;
  LAYER M2 ;
        RECT 6.29 7.84 6.61 8.12 ;
  LAYER M3 ;
        RECT 6.31 7.98 6.59 18.06 ;
  LAYER M2 ;
        RECT 6.29 17.92 6.61 18.2 ;
  LAYER M2 ;
        RECT 6.29 7.84 6.61 8.12 ;
  LAYER M3 ;
        RECT 6.31 7.82 6.59 8.14 ;
  LAYER M2 ;
        RECT 6.29 17.92 6.61 18.2 ;
  LAYER M3 ;
        RECT 6.31 17.9 6.59 18.22 ;
  LAYER M2 ;
        RECT 6.29 7.84 6.61 8.12 ;
  LAYER M3 ;
        RECT 6.31 7.82 6.59 8.14 ;
  LAYER M2 ;
        RECT 6.29 17.92 6.61 18.2 ;
  LAYER M3 ;
        RECT 6.31 17.9 6.59 18.22 ;
  LAYER M2 ;
        RECT 1.12 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 1.12 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 6.28 2.8 9.2 3.08 ;
  LAYER M2 ;
        RECT 6.28 12.04 9.2 12.32 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 7.14 4.01 7.98 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M2 ;
        RECT 3.87 7 5.16 7.28 ;
  LAYER M1 ;
        RECT 5.035 2.94 5.285 7.14 ;
  LAYER M2 ;
        RECT 5.16 2.8 6.45 3.08 ;
  LAYER M1 ;
        RECT 5.035 7.14 5.285 12.18 ;
  LAYER M2 ;
        RECT 5.16 12.04 6.45 12.32 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M1 ;
        RECT 5.035 2.855 5.285 3.025 ;
  LAYER M2 ;
        RECT 4.99 2.8 5.33 3.08 ;
  LAYER M1 ;
        RECT 5.035 7.055 5.285 7.225 ;
  LAYER M2 ;
        RECT 4.99 7 5.33 7.28 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M1 ;
        RECT 5.035 2.855 5.285 3.025 ;
  LAYER M2 ;
        RECT 4.99 2.8 5.33 3.08 ;
  LAYER M1 ;
        RECT 5.035 7.055 5.285 7.225 ;
  LAYER M2 ;
        RECT 4.99 7 5.33 7.28 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M1 ;
        RECT 5.035 2.855 5.285 3.025 ;
  LAYER M2 ;
        RECT 4.99 2.8 5.33 3.08 ;
  LAYER M1 ;
        RECT 5.035 7.055 5.285 7.225 ;
  LAYER M2 ;
        RECT 4.99 7 5.33 7.28 ;
  LAYER M1 ;
        RECT 5.035 12.095 5.285 12.265 ;
  LAYER M2 ;
        RECT 4.99 12.04 5.33 12.32 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M1 ;
        RECT 5.035 2.855 5.285 3.025 ;
  LAYER M2 ;
        RECT 4.99 2.8 5.33 3.08 ;
  LAYER M1 ;
        RECT 5.035 7.055 5.285 7.225 ;
  LAYER M2 ;
        RECT 4.99 7 5.33 7.28 ;
  LAYER M1 ;
        RECT 5.035 12.095 5.285 12.265 ;
  LAYER M2 ;
        RECT 4.99 12.04 5.33 12.32 ;
  LAYER M2 ;
        RECT 3.71 7 4.03 7.28 ;
  LAYER M3 ;
        RECT 3.73 6.98 4.01 7.3 ;
  LAYER M2 ;
        RECT 3.71 7.84 4.03 8.12 ;
  LAYER M3 ;
        RECT 3.73 7.82 4.01 8.14 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 11.425 ;
  LAYER M1 ;
        RECT 2.025 11.675 2.275 12.685 ;
  LAYER M1 ;
        RECT 2.025 13.775 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.455 7.895 2.705 11.425 ;
  LAYER M1 ;
        RECT 2.885 7.895 3.135 11.425 ;
  LAYER M1 ;
        RECT 2.885 11.675 3.135 12.685 ;
  LAYER M1 ;
        RECT 2.885 13.775 3.135 14.785 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 1.12 14.14 4.04 14.42 ;
  LAYER M2 ;
        RECT 1.12 7.84 4.04 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 4.04 12.32 ;
  LAYER M3 ;
        RECT 2.87 8.24 3.15 14.44 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 11.425 ;
  LAYER M1 ;
        RECT 8.905 11.675 9.155 12.685 ;
  LAYER M1 ;
        RECT 8.905 13.775 9.155 14.785 ;
  LAYER M1 ;
        RECT 9.335 7.895 9.585 11.425 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 14.785 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 11.425 ;
  LAYER M1 ;
        RECT 7.185 11.675 7.435 12.685 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M2 ;
        RECT 5.85 8.26 9.63 8.54 ;
  LAYER M2 ;
        RECT 6.28 14.14 9.2 14.42 ;
  LAYER M2 ;
        RECT 6.28 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 6.28 12.04 9.2 12.32 ;
  LAYER M3 ;
        RECT 7.17 8.24 7.45 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 2.025 3.695 2.275 7.225 ;
  LAYER M1 ;
        RECT 2.025 2.435 2.275 3.445 ;
  LAYER M1 ;
        RECT 2.025 0.335 2.275 1.345 ;
  LAYER M1 ;
        RECT 2.455 3.695 2.705 7.225 ;
  LAYER M1 ;
        RECT 2.885 3.695 3.135 7.225 ;
  LAYER M1 ;
        RECT 2.885 2.435 3.135 3.445 ;
  LAYER M1 ;
        RECT 2.885 0.335 3.135 1.345 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M2 ;
        RECT 0.69 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 1.12 0.7 4.04 0.98 ;
  LAYER M2 ;
        RECT 1.12 7 4.04 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 4.04 3.08 ;
  LAYER M3 ;
        RECT 2.87 0.68 3.15 6.88 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M1 ;
        RECT 8.045 3.695 8.295 7.225 ;
  LAYER M1 ;
        RECT 8.045 2.435 8.295 3.445 ;
  LAYER M1 ;
        RECT 8.045 0.335 8.295 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M2 ;
        RECT 5.85 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 6.28 0.7 9.2 0.98 ;
  LAYER M2 ;
        RECT 6.28 7 9.2 7.28 ;
  LAYER M2 ;
        RECT 6.28 2.8 9.2 3.08 ;
  LAYER M3 ;
        RECT 7.17 0.68 7.45 6.88 ;
  LAYER M1 ;
        RECT 6.325 23.015 6.575 26.545 ;
  LAYER M1 ;
        RECT 6.325 26.795 6.575 27.805 ;
  LAYER M1 ;
        RECT 6.325 28.895 6.575 29.905 ;
  LAYER M1 ;
        RECT 6.755 23.015 7.005 26.545 ;
  LAYER M1 ;
        RECT 5.895 23.015 6.145 26.545 ;
  LAYER M1 ;
        RECT 5.465 23.015 5.715 26.545 ;
  LAYER M1 ;
        RECT 5.465 26.795 5.715 27.805 ;
  LAYER M1 ;
        RECT 5.465 28.895 5.715 29.905 ;
  LAYER M1 ;
        RECT 5.035 23.015 5.285 26.545 ;
  LAYER M1 ;
        RECT 4.605 23.015 4.855 26.545 ;
  LAYER M1 ;
        RECT 4.605 26.795 4.855 27.805 ;
  LAYER M1 ;
        RECT 4.605 28.895 4.855 29.905 ;
  LAYER M1 ;
        RECT 4.175 23.015 4.425 26.545 ;
  LAYER M1 ;
        RECT 3.745 23.015 3.995 26.545 ;
  LAYER M1 ;
        RECT 3.745 26.795 3.995 27.805 ;
  LAYER M1 ;
        RECT 3.745 28.895 3.995 29.905 ;
  LAYER M1 ;
        RECT 3.315 23.015 3.565 26.545 ;
  LAYER M2 ;
        RECT 3.27 23.38 7.05 23.66 ;
  LAYER M2 ;
        RECT 3.7 29.26 6.62 29.54 ;
  LAYER M2 ;
        RECT 3.7 22.96 6.62 23.24 ;
  LAYER M2 ;
        RECT 3.7 27.16 6.62 27.44 ;
  LAYER M3 ;
        RECT 4.59 23.36 4.87 29.56 ;
  LAYER M1 ;
        RECT 6.325 18.815 6.575 22.345 ;
  LAYER M1 ;
        RECT 6.325 17.555 6.575 18.565 ;
  LAYER M1 ;
        RECT 6.325 15.455 6.575 16.465 ;
  LAYER M1 ;
        RECT 6.755 18.815 7.005 22.345 ;
  LAYER M1 ;
        RECT 5.895 18.815 6.145 22.345 ;
  LAYER M1 ;
        RECT 5.465 18.815 5.715 22.345 ;
  LAYER M1 ;
        RECT 5.465 17.555 5.715 18.565 ;
  LAYER M1 ;
        RECT 5.465 15.455 5.715 16.465 ;
  LAYER M1 ;
        RECT 5.035 18.815 5.285 22.345 ;
  LAYER M1 ;
        RECT 4.605 18.815 4.855 22.345 ;
  LAYER M1 ;
        RECT 4.605 17.555 4.855 18.565 ;
  LAYER M1 ;
        RECT 4.605 15.455 4.855 16.465 ;
  LAYER M1 ;
        RECT 4.175 18.815 4.425 22.345 ;
  LAYER M1 ;
        RECT 3.745 18.815 3.995 22.345 ;
  LAYER M1 ;
        RECT 3.745 17.555 3.995 18.565 ;
  LAYER M1 ;
        RECT 3.745 15.455 3.995 16.465 ;
  LAYER M1 ;
        RECT 3.315 18.815 3.565 22.345 ;
  LAYER M2 ;
        RECT 3.27 21.7 7.05 21.98 ;
  LAYER M2 ;
        RECT 3.7 15.82 6.62 16.1 ;
  LAYER M2 ;
        RECT 3.7 22.12 6.62 22.4 ;
  LAYER M2 ;
        RECT 3.7 17.92 6.62 18.2 ;
  LAYER M3 ;
        RECT 4.59 15.8 4.87 22 ;
  END 
END RINGOSCILLATOR
