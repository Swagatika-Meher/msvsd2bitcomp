* SPICE3 file created from FUNCTION_0.ext - technology: sky130A

.subckt NMOS_S_21929916_X1_Y1_1677566905_1677566908 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_230_483# a_200_252# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt PMOS_S_95864420_X1_Y1_1677566906_1677566908 a_230_462# a_200_252# w_0_0# VSUBS
X0 a_230_462# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.94e+11p pd=2.66e+06u as=5.565e+11p ps=5.26e+06u w=1.05e+06u l=150000u
X1 w_0_0# a_200_252# a_230_462# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
C0 a_200_252# w_0_0# 0.77fF
C1 a_200_252# a_230_462# 0.11fF
C2 a_230_462# w_0_0# 0.78fF
C3 a_230_462# VSUBS -0.04fF
C4 a_200_252# VSUBS 0.08fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt INV_33643809_0_0_1677566908 m1_312_1400# li_405_571# PMOS_S_95864420_X1_Y1_1677566906_1677566908_0/w_0_0#
+ VSUBS
XNMOS_S_21929916_X1_Y1_1677566905_1677566908_0 li_405_571# m1_312_1400# VSUBS NMOS_S_21929916_X1_Y1_1677566905_1677566908
XPMOS_S_95864420_X1_Y1_1677566906_1677566908_0 m1_312_1400# li_405_571# PMOS_S_95864420_X1_Y1_1677566906_1677566908_0/w_0_0#
+ VSUBS PMOS_S_95864420_X1_Y1_1677566906_1677566908
C0 m1_312_1400# PMOS_S_95864420_X1_Y1_1677566906_1677566908_0/w_0_0# 0.01fF
C1 li_405_571# m1_312_1400# 0.09fF
C2 li_405_571# PMOS_S_95864420_X1_Y1_1677566906_1677566908_0/w_0_0# 0.34fF
C3 m1_312_1400# VSUBS 0.69fF
C4 li_405_571# VSUBS 1.50fF
C5 PMOS_S_95864420_X1_Y1_1677566906_1677566908_0/w_0_0# VSUBS 3.02fF
.ends

.subckt NMOS_S_21929916_X1_Y1_1677566910 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_200_252# a_230_483# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt PMOS_S_95864420_X1_Y1_1677566911 a_230_462# a_200_252# w_0_0# VSUBS
X0 a_230_462# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.94e+11p pd=2.66e+06u as=5.565e+11p ps=5.26e+06u w=1.05e+06u l=150000u
X1 w_0_0# a_200_252# a_230_462# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
C0 a_230_462# a_200_252# 0.11fF
C1 w_0_0# a_200_252# 0.77fF
C2 a_230_462# w_0_0# 0.78fF
C3 a_230_462# VSUBS -0.04fF
C4 a_200_252# VSUBS 0.08fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt DP_PMOS_65570828_X1_Y1_1677566909 a_372_252# a_230_462# a_200_252# a_402_462#
+ w_0_0# VSUBS
X0 w_0_0# a_372_252# a_402_462# w_0_0# sky130_fd_pr__pfet_01v8 ad=8.505e+11p pd=7.92e+06u as=2.94e+11p ps=2.66e+06u w=1.05e+06u l=150000u
X1 a_230_462# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.94e+11p pd=2.66e+06u as=0p ps=0u w=1.05e+06u l=150000u
X2 w_0_0# a_200_252# a_230_462# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
X3 a_402_462# a_372_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.05e+06u l=150000u
C0 a_372_252# a_200_252# 0.25fF
C1 a_200_252# a_402_462# 0.01fF
C2 a_372_252# a_402_462# 0.11fF
C3 w_0_0# a_200_252# 0.65fF
C4 a_372_252# w_0_0# 0.66fF
C5 a_230_462# a_200_252# 0.12fF
C6 w_0_0# a_402_462# 0.91fF
C7 a_230_462# a_402_462# 0.06fF
C8 a_230_462# w_0_0# 0.72fF
C9 a_402_462# VSUBS -0.06fF
C10 a_230_462# VSUBS -0.11fF
C11 a_372_252# VSUBS 0.05fF
C12 a_200_252# VSUBS 0.01fF
C13 w_0_0# VSUBS 3.45fF
.ends

.subckt FUNCTION_0
XINV_33643809_0_0_1677566908_0 FN E VDD GND INV_33643809_0_0_1677566908
XNMOS_S_21929916_X1_Y1_1677566910_0 li_2469_571# FN GND NMOS_S_21929916_X1_Y1_1677566910
XNMOS_S_21929916_X1_Y1_1677566910_1 m1_1430_896# FN GND NMOS_S_21929916_X1_Y1_1677566910
XNMOS_S_21929916_X1_Y1_1677566910_2 F GND GND NMOS_S_21929916_X1_Y1_1677566910
XNMOS_S_21929916_X1_Y1_1677566910_3 D GND GND NMOS_S_21929916_X1_Y1_1677566910
XNMOS_S_21929916_X1_Y1_1677566910_4 B GND GND NMOS_S_21929916_X1_Y1_1677566910
XPMOS_S_95864420_X1_Y1_1677566911_0 FN F VDD GND PMOS_S_95864420_X1_Y1_1677566911
XPMOS_S_95864420_X1_Y1_1677566911_1 VDD D VDD GND PMOS_S_95864420_X1_Y1_1677566911
XPMOS_S_95864420_X1_Y1_1677566911_2 VDD li_2469_571# VDD GND PMOS_S_95864420_X1_Y1_1677566911
XDP_PMOS_65570828_X1_Y1_1677566909_0 B VDD m1_1430_896# VDD VDD GND DP_PMOS_65570828_X1_Y1_1677566909
C0 VDD F 0.62fF
C1 m1_1430_896# D 0.15fF
C2 B m1_1430_896# 0.03fF
C3 A FN -0.00fF
C4 VDD D 0.75fF
C5 B VDD 1.08fF
C6 li_2469_571# D 0.05fF
C7 F FN 0.20fF
C8 B li_2469_571# 0.14fF
C9 A F -0.01fF
C10 FN D 0.01fF
C11 A D 0.15fF
C12 B A -0.02fF
C13 F D 0.01fF
C14 B F 0.00fF
C15 VDD C 0.78fF
C16 VDD E 0.06fF
C17 B D 0.00fF
C18 VDD m1_1430_896# 0.10fF
C19 FN C -0.00fF
C20 A C 0.00fF
C21 FN E 0.03fF
C22 m1_1430_896# li_2469_571# 0.00fF
C23 A E 0.00fF
C24 VDD li_2469_571# 0.04fF
C25 m1_1430_896# FN 0.00fF
C26 F E 0.03fF
C27 VDD FN 1.61fF
C28 A VDD 1.01fF
C29 C D 0.01fF
C30 E D 0.01fF
C31 B C 0.13fF
C32 FN li_2469_571# -0.00fF
C33 m1_1430_896# F 0.07fF
C34 C GND 0.19fF **FLOATING
C35 A GND 0.11fF **FLOATING
C36 B GND 1.70fF
C37 D GND 1.93fF
C38 F GND 0.71fF
C39 m1_1430_896# GND 1.45fF
C40 li_2469_571# GND 1.77fF
C41 FN GND 1.59fF
C42 E GND 1.19fF
C43 VDD GND 14.04fF
.ends

