* NGSPICE file created from function_post.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
C0 a_n73_n100# a_n33_n188# 0.03fF
C1 a_15_n100# a_n73_n100# 0.16fF
C2 a_15_n100# a_n33_n188# 0.03fF
C3 a_15_n100# a_n175_n274# 0.08fF
C4 a_n73_n100# a_n175_n274# 0.11fF
C5 a_n33_n188# a_n175_n274# 0.30fF
.ends

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
C0 a_15_n100# a_n33_n197# 0.03fF
C1 a_n33_n197# w_n211_n319# 0.26fF
C2 a_n73_n100# a_n33_n197# 0.03fF
C3 a_15_n100# w_n211_n319# 0.06fF
C4 a_15_n100# a_n73_n100# 0.16fF
C5 a_n73_n100# w_n211_n319# 0.09fF
C6 a_15_n100# VSUBS 0.02fF
C7 a_n73_n100# VSUBS 0.02fF
C8 a_n33_n197# VSUBS 0.05fF
C9 w_n211_n319# VSUBS 1.07fF
.ends

.subckt function_post VDD A B D C F E Fn Gnd
XXM12 m1_n4122_n2248# F Gnd VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM1 VDD m1_n6798_n26# XM1/w_n211_n319# A VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM2 m1_n638_22# VDD XM2/w_n211_n319# B VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM3 m1_n6798_n26# m1_n5500_n14# XM3/w_n211_n319# C VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM4 m1_n5500_n14# m1_n638_22# XM4/w_n211_n319# D VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM5 m1_n5500_n14# Fn XM5/w_n211_n319# E VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM6 Fn m1_n5500_n14# XM6/w_n211_n319# F VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM7 Fn A m1_n7132_n2270# VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM9 Fn E m1_n4122_n2248# VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM8 m1_n7132_n2270# C Fn VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM10 m1_n7132_n2270# B Gnd VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM11 Gnd D m1_n7132_n2270# VSUBS sky130_fd_pr__nfet_01v8_648S5X
C0 XM2/w_n211_n319# B 0.10fF
C1 XM6/w_n211_n319# D 0.00fF
C2 XM4/w_n211_n319# m1_n5500_n14# 0.07fF
C3 VDD C 0.01fF
C4 m1_n5500_n14# XM3/w_n211_n319# 0.08fF
C5 Fn m1_n7132_n2270# 0.10fF
C6 m1_n7132_n2270# F 0.00fF
C7 Fn E 0.29fF
C8 F E 0.01fF
C9 VDD XM5/w_n211_n319# 0.04fF
C10 XM1/w_n211_n319# A 0.12fF
C11 A Fn 0.17fF
C12 VDD m1_n5500_n14# 1.48fF
C13 C m1_n7132_n2270# 0.01fF
C14 C E 0.07fF
C15 XM1/w_n211_n319# m1_n6798_n26# 0.08fF
C16 Fn m1_n6798_n26# 0.00fF
C17 m1_n638_22# B 0.01fF
C18 VDD XM4/w_n211_n319# 0.03fF
C19 C A 0.07fF
C20 VDD XM3/w_n211_n319# 0.04fF
C21 XM5/w_n211_n319# E 0.10fF
C22 XM2/w_n211_n319# D 0.00fF
C23 C m1_n6798_n26# 0.01fF
C24 m1_n5500_n14# E 0.01fF
C25 XM6/w_n211_n319# Fn 0.09fF
C26 XM6/w_n211_n319# F 0.05fF
C27 A m1_n5500_n14# 0.00fF
C28 XM3/w_n211_n319# E 0.00fF
C29 m1_n5500_n14# m1_n6798_n26# 0.00fF
C30 A XM3/w_n211_n319# 0.00fF
C31 XM6/w_n211_n319# XM5/w_n211_n319# 0.01fF
C32 m1_n638_22# D 0.01fF
C33 Gnd m1_n7132_n2270# 0.83fF
C34 D F 0.01fF
C35 XM4/w_n211_n319# B 0.00fF
C36 XM3/w_n211_n319# m1_n6798_n26# 0.07fF
C37 VDD E 0.01fF
C38 XM6/w_n211_n319# m1_n5500_n14# 0.12fF
C39 VDD A 0.03fF
C40 m1_n638_22# XM2/w_n211_n319# 0.07fF
C41 XM6/w_n211_n319# XM4/w_n211_n319# 0.01fF
C42 Gnd B 0.02fF
C43 VDD m1_n6798_n26# 0.06fF
C44 VDD B 0.02fF
C45 m1_n7132_n2270# E 0.00fF
C46 Fn m1_n4122_n2248# 0.04fF
C47 F m1_n4122_n2248# 0.00fF
C48 A m1_n7132_n2270# 0.02fF
C49 m1_n5500_n14# D 0.01fF
C50 VDD XM6/w_n211_n319# 0.04fF
C51 C m1_n4122_n2248# 0.00fF
C52 XM4/w_n211_n319# D 0.10fF
C53 XM1/w_n211_n319# Fn 0.00fF
C54 m1_n7132_n2270# B 0.00fF
C55 m1_n6798_n26# E 0.00fF
C56 Fn F 0.04fF
C57 A m1_n6798_n26# 0.01fF
C58 XM4/w_n211_n319# XM2/w_n211_n319# 0.01fF
C59 XM1/w_n211_n319# C 0.00fF
C60 C Fn 0.20fF
C61 XM6/w_n211_n319# E 0.00fF
C62 Gnd D 0.02fF
C63 VDD D 0.01fF
C64 Fn XM5/w_n211_n319# 0.08fF
C65 XM5/w_n211_n319# F 0.00fF
C66 XM1/w_n211_n319# m1_n5500_n14# 0.00fF
C67 VDD XM2/w_n211_n319# 0.11fF
C68 m1_n638_22# m1_n5500_n14# 0.00fF
C69 m1_n5500_n14# Fn 0.07fF
C70 m1_n5500_n14# F 0.01fF
C71 C XM5/w_n211_n319# 0.00fF
C72 m1_n7132_n2270# D 0.01fF
C73 m1_n638_22# XM4/w_n211_n319# 0.07fF
C74 Gnd m1_n4122_n2248# 0.00fF
C75 XM4/w_n211_n319# F 0.00fF
C76 XM1/w_n211_n319# XM3/w_n211_n319# 0.01fF
C77 XM3/w_n211_n319# Fn 0.01fF
C78 C m1_n5500_n14# 0.01fF
C79 m1_n5500_n14# XM5/w_n211_n319# 0.09fF
C80 C XM3/w_n211_n319# 0.14fF
C81 D B 0.06fF
C82 Gnd F 0.01fF
C83 VDD XM1/w_n211_n319# 0.11fF
C84 VDD m1_n638_22# 0.08fF
C85 VDD Fn 0.08fF
C86 VDD F 0.01fF
C87 m1_n7132_n2270# m1_n4122_n2248# 0.00fF
C88 E m1_n4122_n2248# 0.00fF
C89 XM3/w_n211_n319# XM5/w_n211_n319# 0.01fF
C90 D VSUBS 1.06fF
C91 B VSUBS 1.06fF
C92 F VSUBS 1.13fF
C93 E VSUBS 1.00fF
C94 C VSUBS 0.91fF
C95 A VSUBS 1.12fF
C96 m1_n4122_n2248# VSUBS 0.66fF
C97 m1_n7132_n2270# VSUBS 2.52fF
C98 Fn VSUBS 3.63fF
C99 XM6/w_n211_n319# VSUBS 1.07fF
C100 XM5/w_n211_n319# VSUBS 1.07fF
C101 m1_n638_22# VSUBS -0.27fF
C102 XM4/w_n211_n319# VSUBS 1.07fF
C103 m1_n5500_n14# VSUBS 1.43fF
C104 XM3/w_n211_n319# VSUBS 1.07fF
C105 XM2/w_n211_n319# VSUBS 1.07fF
C106 m1_n6798_n26# VSUBS 0.00fF
C107 VDD VSUBS 0.53fF
C108 XM1/w_n211_n319# VSUBS 1.07fF
C109 Gnd VSUBS 2.79fF
.ends


*========Manually added===========

V1 A GND pulse(0 1.8 0.1n 10p 10p 1n 2n)
.save i(v1)
V2 B GND pulse(0 1.8 0.2n 10p 10p 1n 2n)
.save i(v2)
V3 C GND pulse(0 1.8 0.3n 10p 10p 1n 2n)
.save i(v3)
V4 D GND pulse(0 1.8 0.4n 10p 10p 1n 2n)
.save i(v4)
V5 E GND pulse(0 1.8 0.5n 10p 10p 1n 2n)
.save i(v5)
V6 F GND pulse(0 1.8 0.6n 10p 10p 1n 2n)
.save i(v6)
V7 VDD GND 1.8
.save i(v7)
x1 VDD A B D C F E Fn GND function_post
**** begin user architecture code


.tran 10p 4n
.control
run
plot A+3 B+3 C+3 D+3 E+3 F+3 Fn
.save all
.endc
.end


.lib /home/swagatika/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.save all
.GLOBAL GND
.end


