MACRO FUNCTION
  ORIGIN 0 0 ;
  FOREIGN FUNCTION 0 0 ;
  SIZE 15.48 BY 15.12 ;
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
      LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
      LAYER M2 ;
        RECT 0.27 2.8 0.59 3.08 ;
      LAYER M1 ;
        RECT 0.305 2.94 0.555 12.18 ;
      LAYER M2 ;
        RECT 0.27 12.04 0.59 12.32 ;
    END
  END E
  PIN FN
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
      LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
      LAYER M2 ;
        RECT 0.7 7 1.02 7.28 ;
      LAYER M3 ;
        RECT 0.72 7.14 1 7.98 ;
      LAYER M2 ;
        RECT 0.7 7.84 1.02 8.12 ;
      LAYER M2 ;
        RECT 2.84 14.56 4.04 14.84 ;
      LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
      LAYER M2 ;
        RECT 11.44 14.56 12.64 14.84 ;
      LAYER M2 ;
        RECT 1.29 7.84 3.01 8.12 ;
      LAYER M1 ;
        RECT 2.885 7.98 3.135 14.7 ;
      LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
      LAYER M2 ;
        RECT 3.87 14.56 6.45 14.84 ;
      LAYER M2 ;
        RECT 7.15 14.56 7.47 14.84 ;
      LAYER M1 ;
        RECT 7.185 14.7 7.435 15.12 ;
      LAYER M2 ;
        RECT 7.31 14.98 9.89 15.26 ;
      LAYER M1 ;
        RECT 9.765 14.7 10.015 15.12 ;
      LAYER M2 ;
        RECT 9.89 14.56 11.61 14.84 ;
    END
  END FN
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.86 4.48 10.06 4.76 ;
      LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
      LAYER M2 ;
        RECT 7.31 4.48 9.03 4.76 ;
      LAYER M3 ;
        RECT 7.17 4.62 7.45 10.5 ;
      LAYER M2 ;
        RECT 7.15 10.36 7.47 10.64 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 9.72 4.9 10.92 5.18 ;
      LAYER M2 ;
        RECT 13.16 10.36 14.36 10.64 ;
      LAYER M2 ;
        RECT 10.75 4.9 13.33 5.18 ;
      LAYER M3 ;
        RECT 13.19 5.04 13.47 10.5 ;
      LAYER M2 ;
        RECT 13.17 10.36 13.49 10.64 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 11.04 1.1 11.32 6.88 ;
    END
  END VDD
  PIN GND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
      LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
      LAYER M3 ;
        RECT 14.48 8.24 14.76 14.44 ;
      LAYER M3 ;
        RECT 4.16 6.115 4.44 6.485 ;
      LAYER M2 ;
        RECT 4.3 6.16 9.46 6.44 ;
      LAYER M3 ;
        RECT 9.32 6.3 9.6 8.4 ;
      LAYER M3 ;
        RECT 9.32 8.635 9.6 9.005 ;
      LAYER M2 ;
        RECT 9.46 8.68 14.62 8.96 ;
      LAYER M3 ;
        RECT 14.48 8.635 14.76 9.005 ;
    END
  END GND
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 7.14 2.8 8.34 3.08 ;
      LAYER M2 ;
        RECT 8 10.36 9.2 10.64 ;
      LAYER M2 ;
        RECT 8.01 2.8 8.33 3.08 ;
      LAYER M1 ;
        RECT 8.045 2.94 8.295 10.5 ;
      LAYER M2 ;
        RECT 8.01 10.36 8.33 10.64 ;
    END
  END D
  PIN F
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 2.84 4.48 4.04 4.76 ;
      LAYER M2 ;
        RECT 2.84 10.36 4.04 10.64 ;
      LAYER M2 ;
        RECT 3.28 4.48 3.6 4.76 ;
      LAYER M3 ;
        RECT 3.3 4.62 3.58 10.5 ;
      LAYER M2 ;
        RECT 3.28 10.36 3.6 10.64 ;
    END
  END F
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 12.3 2.8 13.5 3.08 ;
      LAYER M2 ;
        RECT 11.44 10.36 12.64 10.64 ;
      LAYER M2 ;
        RECT 12.31 2.8 12.63 3.08 ;
      LAYER M1 ;
        RECT 12.345 2.94 12.595 10.5 ;
      LAYER M2 ;
        RECT 12.31 10.36 12.63 10.64 ;
    END
  END C
  OBS 
  LAYER M2 ;
        RECT 2.84 0.28 4.04 0.56 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M2 ;
        RECT 1.72 0.28 3.01 0.56 ;
  LAYER M3 ;
        RECT 1.58 0.42 1.86 0.84 ;
  LAYER M2 ;
        RECT 1.56 0.28 1.88 0.56 ;
  LAYER M3 ;
        RECT 1.58 0.26 1.86 0.58 ;
  LAYER M2 ;
        RECT 1.56 0.28 1.88 0.56 ;
  LAYER M3 ;
        RECT 1.58 0.26 1.86 0.58 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
  LAYER M2 ;
        RECT 7.14 7 8.34 7.28 ;
  LAYER M2 ;
        RECT 12.3 7 13.5 7.28 ;
  LAYER M3 ;
        RECT 1.58 9.055 1.86 9.425 ;
  LAYER M2 ;
        RECT 1.72 9.1 4.3 9.38 ;
  LAYER M3 ;
        RECT 4.16 9.055 4.44 9.425 ;
  LAYER M3 ;
        RECT 4.16 7.56 4.44 8.4 ;
  LAYER M2 ;
        RECT 4.3 7.42 6.45 7.7 ;
  LAYER M1 ;
        RECT 6.325 7.14 6.575 7.56 ;
  LAYER M2 ;
        RECT 6.45 7 7.31 7.28 ;
  LAYER M2 ;
        RECT 8.17 7 12.47 7.28 ;
  LAYER M2 ;
        RECT 1.56 9.1 1.88 9.38 ;
  LAYER M3 ;
        RECT 1.58 9.08 1.86 9.4 ;
  LAYER M2 ;
        RECT 4.14 9.1 4.46 9.38 ;
  LAYER M3 ;
        RECT 4.16 9.08 4.44 9.4 ;
  LAYER M2 ;
        RECT 1.56 9.1 1.88 9.38 ;
  LAYER M3 ;
        RECT 1.58 9.08 1.86 9.4 ;
  LAYER M2 ;
        RECT 4.14 9.1 4.46 9.38 ;
  LAYER M3 ;
        RECT 4.16 9.08 4.44 9.4 ;
  LAYER M1 ;
        RECT 6.325 7.055 6.575 7.225 ;
  LAYER M2 ;
        RECT 6.28 7 6.62 7.28 ;
  LAYER M1 ;
        RECT 6.325 7.475 6.575 7.645 ;
  LAYER M2 ;
        RECT 6.28 7.42 6.62 7.7 ;
  LAYER M2 ;
        RECT 1.56 9.1 1.88 9.38 ;
  LAYER M3 ;
        RECT 1.58 9.08 1.86 9.4 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M2 ;
        RECT 4.14 9.1 4.46 9.38 ;
  LAYER M3 ;
        RECT 4.16 9.08 4.44 9.4 ;
  LAYER M1 ;
        RECT 6.325 7.055 6.575 7.225 ;
  LAYER M2 ;
        RECT 6.28 7 6.62 7.28 ;
  LAYER M1 ;
        RECT 6.325 7.475 6.575 7.645 ;
  LAYER M2 ;
        RECT 6.28 7.42 6.62 7.7 ;
  LAYER M2 ;
        RECT 1.56 9.1 1.88 9.38 ;
  LAYER M3 ;
        RECT 1.58 9.08 1.86 9.4 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M2 ;
        RECT 4.14 9.1 4.46 9.38 ;
  LAYER M3 ;
        RECT 4.16 9.08 4.44 9.4 ;
  LAYER M1 ;
        RECT 6.325 7.055 6.575 7.225 ;
  LAYER M2 ;
        RECT 6.28 7 6.62 7.28 ;
  LAYER M1 ;
        RECT 6.325 7.475 6.575 7.645 ;
  LAYER M2 ;
        RECT 6.28 7.42 6.62 7.7 ;
  LAYER M2 ;
        RECT 1.56 9.1 1.88 9.38 ;
  LAYER M3 ;
        RECT 1.58 9.08 1.86 9.4 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M2 ;
        RECT 4.14 9.1 4.46 9.38 ;
  LAYER M3 ;
        RECT 4.16 9.08 4.44 9.4 ;
  LAYER M1 ;
        RECT 6.325 7.055 6.575 7.225 ;
  LAYER M2 ;
        RECT 6.28 7 6.62 7.28 ;
  LAYER M1 ;
        RECT 6.325 7.475 6.575 7.645 ;
  LAYER M2 ;
        RECT 6.28 7.42 6.62 7.7 ;
  LAYER M2 ;
        RECT 1.56 9.1 1.88 9.38 ;
  LAYER M3 ;
        RECT 1.58 9.08 1.86 9.4 ;
  LAYER M2 ;
        RECT 4.14 7.42 4.46 7.7 ;
  LAYER M3 ;
        RECT 4.16 7.4 4.44 7.72 ;
  LAYER M2 ;
        RECT 4.14 9.1 4.46 9.38 ;
  LAYER M3 ;
        RECT 4.16 9.08 4.44 9.4 ;
  LAYER M2 ;
        RECT 8.86 0.28 10.06 0.56 ;
  LAYER M3 ;
        RECT 13.62 0.68 13.9 6.88 ;
  LAYER M2 ;
        RECT 9.89 0.28 13.76 0.56 ;
  LAYER M3 ;
        RECT 13.62 0.42 13.9 0.84 ;
  LAYER M2 ;
        RECT 13.6 0.28 13.92 0.56 ;
  LAYER M3 ;
        RECT 13.62 0.26 13.9 0.58 ;
  LAYER M2 ;
        RECT 13.6 0.28 13.92 0.56 ;
  LAYER M3 ;
        RECT 13.62 0.26 13.9 0.58 ;
  LAYER M2 ;
        RECT 9.72 0.7 10.92 0.98 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M2 ;
        RECT 8.6 0.7 9.89 0.98 ;
  LAYER M3 ;
        RECT 8.46 0 8.74 0.84 ;
  LAYER M2 ;
        RECT 8.17 -0.14 8.6 0.14 ;
  LAYER M3 ;
        RECT 8.03 0 8.31 0.42 ;
  LAYER M2 ;
        RECT 6.88 0.28 8.17 0.56 ;
  LAYER M3 ;
        RECT 6.74 0.42 7.02 0.84 ;
  LAYER M2 ;
        RECT 6.72 0.28 7.04 0.56 ;
  LAYER M3 ;
        RECT 6.74 0.26 7.02 0.58 ;
  LAYER M2 ;
        RECT 8.01 -0.14 8.33 0.14 ;
  LAYER M3 ;
        RECT 8.03 -0.16 8.31 0.16 ;
  LAYER M2 ;
        RECT 8.01 0.28 8.33 0.56 ;
  LAYER M3 ;
        RECT 8.03 0.26 8.31 0.58 ;
  LAYER M2 ;
        RECT 8.44 -0.14 8.76 0.14 ;
  LAYER M3 ;
        RECT 8.46 -0.16 8.74 0.16 ;
  LAYER M2 ;
        RECT 8.44 0.7 8.76 0.98 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 1 ;
  LAYER M2 ;
        RECT 6.72 0.28 7.04 0.56 ;
  LAYER M3 ;
        RECT 6.74 0.26 7.02 0.58 ;
  LAYER M2 ;
        RECT 8.01 -0.14 8.33 0.14 ;
  LAYER M3 ;
        RECT 8.03 -0.16 8.31 0.16 ;
  LAYER M2 ;
        RECT 8.01 0.28 8.33 0.56 ;
  LAYER M3 ;
        RECT 8.03 0.26 8.31 0.58 ;
  LAYER M2 ;
        RECT 8.44 -0.14 8.76 0.14 ;
  LAYER M3 ;
        RECT 8.46 -0.16 8.74 0.16 ;
  LAYER M2 ;
        RECT 8.44 0.7 8.76 0.98 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 1 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
  LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
  LAYER M2 ;
        RECT 8 14.56 9.2 14.84 ;
  LAYER M2 ;
        RECT 13.16 14.56 14.36 14.84 ;
  LAYER M3 ;
        RECT 5.88 12.835 6.16 13.205 ;
  LAYER M2 ;
        RECT 6.02 12.88 11.18 13.16 ;
  LAYER M3 ;
        RECT 11.04 12.835 11.32 13.205 ;
  LAYER M2 ;
        RECT 8.87 12.88 9.19 13.16 ;
  LAYER M3 ;
        RECT 8.89 13.02 9.17 14.7 ;
  LAYER M2 ;
        RECT 8.87 14.56 9.19 14.84 ;
  LAYER M3 ;
        RECT 11.04 13.675 11.32 14.045 ;
  LAYER M2 ;
        RECT 11.18 13.72 13.33 14 ;
  LAYER M1 ;
        RECT 13.205 13.86 13.455 14.7 ;
  LAYER M2 ;
        RECT 13.17 14.56 13.49 14.84 ;
  LAYER M2 ;
        RECT 5.86 12.88 6.18 13.16 ;
  LAYER M3 ;
        RECT 5.88 12.86 6.16 13.18 ;
  LAYER M2 ;
        RECT 11.02 12.88 11.34 13.16 ;
  LAYER M3 ;
        RECT 11.04 12.86 11.32 13.18 ;
  LAYER M2 ;
        RECT 5.86 12.88 6.18 13.16 ;
  LAYER M3 ;
        RECT 5.88 12.86 6.16 13.18 ;
  LAYER M2 ;
        RECT 11.02 12.88 11.34 13.16 ;
  LAYER M3 ;
        RECT 11.04 12.86 11.32 13.18 ;
  LAYER M2 ;
        RECT 5.86 12.88 6.18 13.16 ;
  LAYER M3 ;
        RECT 5.88 12.86 6.16 13.18 ;
  LAYER M2 ;
        RECT 8.87 12.88 9.19 13.16 ;
  LAYER M3 ;
        RECT 8.89 12.86 9.17 13.18 ;
  LAYER M2 ;
        RECT 8.87 14.56 9.19 14.84 ;
  LAYER M3 ;
        RECT 8.89 14.54 9.17 14.86 ;
  LAYER M2 ;
        RECT 11.02 12.88 11.34 13.16 ;
  LAYER M3 ;
        RECT 11.04 12.86 11.32 13.18 ;
  LAYER M2 ;
        RECT 5.86 12.88 6.18 13.16 ;
  LAYER M3 ;
        RECT 5.88 12.86 6.16 13.18 ;
  LAYER M2 ;
        RECT 8.87 12.88 9.19 13.16 ;
  LAYER M3 ;
        RECT 8.89 12.86 9.17 13.18 ;
  LAYER M2 ;
        RECT 8.87 14.56 9.19 14.84 ;
  LAYER M3 ;
        RECT 8.89 14.54 9.17 14.86 ;
  LAYER M2 ;
        RECT 11.02 12.88 11.34 13.16 ;
  LAYER M3 ;
        RECT 11.04 12.86 11.32 13.18 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 13.945 ;
  LAYER M2 ;
        RECT 13.16 13.72 13.5 14 ;
  LAYER M1 ;
        RECT 13.205 14.615 13.455 14.785 ;
  LAYER M2 ;
        RECT 13.16 14.56 13.5 14.84 ;
  LAYER M2 ;
        RECT 5.86 12.88 6.18 13.16 ;
  LAYER M3 ;
        RECT 5.88 12.86 6.16 13.18 ;
  LAYER M2 ;
        RECT 8.87 12.88 9.19 13.16 ;
  LAYER M3 ;
        RECT 8.89 12.86 9.17 13.18 ;
  LAYER M2 ;
        RECT 8.87 14.56 9.19 14.84 ;
  LAYER M3 ;
        RECT 8.89 14.54 9.17 14.86 ;
  LAYER M2 ;
        RECT 11.02 12.88 11.34 13.16 ;
  LAYER M3 ;
        RECT 11.04 12.86 11.32 13.18 ;
  LAYER M2 ;
        RECT 11.02 13.72 11.34 14 ;
  LAYER M3 ;
        RECT 11.04 13.7 11.32 14.02 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 13.945 ;
  LAYER M2 ;
        RECT 13.16 13.72 13.5 14 ;
  LAYER M1 ;
        RECT 13.205 14.615 13.455 14.785 ;
  LAYER M2 ;
        RECT 13.16 14.56 13.5 14.84 ;
  LAYER M2 ;
        RECT 5.86 12.88 6.18 13.16 ;
  LAYER M3 ;
        RECT 5.88 12.86 6.16 13.18 ;
  LAYER M2 ;
        RECT 8.87 12.88 9.19 13.16 ;
  LAYER M3 ;
        RECT 8.89 12.86 9.17 13.18 ;
  LAYER M2 ;
        RECT 8.87 14.56 9.19 14.84 ;
  LAYER M3 ;
        RECT 8.89 14.54 9.17 14.86 ;
  LAYER M2 ;
        RECT 11.02 12.88 11.34 13.16 ;
  LAYER M3 ;
        RECT 11.04 12.86 11.32 13.18 ;
  LAYER M2 ;
        RECT 11.02 13.72 11.34 14 ;
  LAYER M3 ;
        RECT 11.04 13.7 11.32 14.02 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 9.765 0.335 10.015 3.865 ;
  LAYER M1 ;
        RECT 9.765 4.115 10.015 5.125 ;
  LAYER M1 ;
        RECT 9.765 6.215 10.015 7.225 ;
  LAYER M1 ;
        RECT 9.335 0.335 9.585 3.865 ;
  LAYER M1 ;
        RECT 10.195 0.335 10.445 3.865 ;
  LAYER M1 ;
        RECT 10.625 0.335 10.875 3.865 ;
  LAYER M1 ;
        RECT 10.625 4.115 10.875 5.125 ;
  LAYER M1 ;
        RECT 10.625 6.215 10.875 7.225 ;
  LAYER M1 ;
        RECT 11.055 0.335 11.305 3.865 ;
  LAYER M2 ;
        RECT 9.72 6.58 11.35 6.86 ;
  LAYER M2 ;
        RECT 9.29 1.12 11.35 1.4 ;
  LAYER M2 ;
        RECT 8.86 0.28 10.06 0.56 ;
  LAYER M2 ;
        RECT 9.72 0.7 10.92 0.98 ;
  LAYER M2 ;
        RECT 8.86 4.48 10.06 4.76 ;
  LAYER M2 ;
        RECT 9.72 4.9 10.92 5.18 ;
  LAYER M3 ;
        RECT 11.04 1.1 11.32 6.88 ;
  LAYER M1 ;
        RECT 14.065 11.255 14.315 14.785 ;
  LAYER M1 ;
        RECT 14.065 9.995 14.315 11.005 ;
  LAYER M1 ;
        RECT 14.065 7.895 14.315 8.905 ;
  LAYER M1 ;
        RECT 13.635 11.255 13.885 14.785 ;
  LAYER M1 ;
        RECT 14.495 11.255 14.745 14.785 ;
  LAYER M2 ;
        RECT 13.59 8.26 14.79 8.54 ;
  LAYER M2 ;
        RECT 13.59 14.14 14.79 14.42 ;
  LAYER M2 ;
        RECT 13.16 14.56 14.36 14.84 ;
  LAYER M2 ;
        RECT 13.16 10.36 14.36 10.64 ;
  LAYER M3 ;
        RECT 14.48 8.24 14.76 14.44 ;
  LAYER M1 ;
        RECT 8.905 11.255 9.155 14.785 ;
  LAYER M1 ;
        RECT 8.905 9.995 9.155 11.005 ;
  LAYER M1 ;
        RECT 8.905 7.895 9.155 8.905 ;
  LAYER M1 ;
        RECT 8.475 11.255 8.725 14.785 ;
  LAYER M1 ;
        RECT 9.335 11.255 9.585 14.785 ;
  LAYER M2 ;
        RECT 8.43 8.26 9.63 8.54 ;
  LAYER M2 ;
        RECT 8.43 14.14 9.63 14.42 ;
  LAYER M2 ;
        RECT 8 14.56 9.2 14.84 ;
  LAYER M2 ;
        RECT 8 10.36 9.2 10.64 ;
  LAYER M3 ;
        RECT 9.32 8.24 9.6 14.44 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 3.865 ;
  LAYER M1 ;
        RECT 3.745 4.115 3.995 5.125 ;
  LAYER M1 ;
        RECT 3.745 6.215 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.315 0.335 3.565 3.865 ;
  LAYER M1 ;
        RECT 4.175 0.335 4.425 3.865 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 2.84 0.28 4.04 0.56 ;
  LAYER M2 ;
        RECT 2.84 4.48 4.04 4.76 ;
  LAYER M3 ;
        RECT 4.16 0.68 4.44 6.88 ;
  LAYER M1 ;
        RECT 6.325 11.255 6.575 14.785 ;
  LAYER M1 ;
        RECT 6.325 9.995 6.575 11.005 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 8.905 ;
  LAYER M1 ;
        RECT 6.755 11.255 7.005 14.785 ;
  LAYER M1 ;
        RECT 5.895 11.255 6.145 14.785 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 6.28 14.56 7.48 14.84 ;
  LAYER M2 ;
        RECT 6.28 10.36 7.48 10.64 ;
  LAYER M3 ;
        RECT 5.88 8.24 6.16 14.44 ;
  LAYER M1 ;
        RECT 11.485 11.255 11.735 14.785 ;
  LAYER M1 ;
        RECT 11.485 9.995 11.735 11.005 ;
  LAYER M1 ;
        RECT 11.485 7.895 11.735 8.905 ;
  LAYER M1 ;
        RECT 11.915 11.255 12.165 14.785 ;
  LAYER M1 ;
        RECT 11.055 11.255 11.305 14.785 ;
  LAYER M2 ;
        RECT 11.01 8.26 12.21 8.54 ;
  LAYER M2 ;
        RECT 11.01 14.14 12.21 14.42 ;
  LAYER M2 ;
        RECT 11.44 14.56 12.64 14.84 ;
  LAYER M2 ;
        RECT 11.44 10.36 12.64 10.64 ;
  LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
  LAYER M1 ;
        RECT 13.205 3.695 13.455 7.225 ;
  LAYER M1 ;
        RECT 13.205 2.435 13.455 3.445 ;
  LAYER M1 ;
        RECT 13.205 0.335 13.455 1.345 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M1 ;
        RECT 13.635 3.695 13.885 7.225 ;
  LAYER M2 ;
        RECT 12.73 0.7 13.93 0.98 ;
  LAYER M2 ;
        RECT 12.73 6.58 13.93 6.86 ;
  LAYER M2 ;
        RECT 12.3 7 13.5 7.28 ;
  LAYER M2 ;
        RECT 12.3 2.8 13.5 3.08 ;
  LAYER M3 ;
        RECT 13.62 0.68 13.9 6.88 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 6.71 0.7 7.91 0.98 ;
  LAYER M2 ;
        RECT 6.71 6.58 7.91 6.86 ;
  LAYER M2 ;
        RECT 7.14 7 8.34 7.28 ;
  LAYER M2 ;
        RECT 7.14 2.8 8.34 3.08 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M1 ;
        RECT 3.745 11.255 3.995 14.785 ;
  LAYER M1 ;
        RECT 3.745 9.995 3.995 11.005 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 8.905 ;
  LAYER M1 ;
        RECT 3.315 11.255 3.565 14.785 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 2.84 14.56 4.04 14.84 ;
  LAYER M2 ;
        RECT 2.84 10.36 4.04 10.64 ;
  LAYER M3 ;
        RECT 4.16 8.24 4.44 14.44 ;
  END 
END FUNCTION
