* SPICE3 file created from flash_adc.ext - technology: sky130A

.subckt flash_adc T_1 T_6 T_7 VIN T_2 T_3 T_4 T_5 Y1 Y2 Y3 VDD GND
X0 T_4 FLASH_ADC_SYM_4_0/a_200_531# VDD VDD sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.41903e+13p ps=4.3592e+08u w=840000u l=150000u
X1 VDD VIN FLASH_ADC_SYM_4_0/a_200_531# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=2.352e+11p ps=2.24e+06u w=840000u l=150000u
X2 VDD FLASH_ADC_SYM_4_0/a_200_531# T_4 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 T_4 FLASH_ADC_SYM_4_0/a_200_531# GND GND sky130_fd_pr__nfet_01v8 ad=4.704e+11p pd=3.92e+06u as=3.09329e+13p ps=3.3716e+08u w=1.68e+06u l=150000u
X4 GND FLASH_ADC_SYM_4_0/a_200_531# T_4 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X5 FLASH_ADC_SYM_4_0/a_200_531# VIN GND GND sky130_fd_pr__nfet_01v8 ad=4.704e+11p pd=3.92e+06u as=0p ps=0u w=1.68e+06u l=150000u
X6 GND VIN FLASH_ADC_SYM_4_0/a_200_531# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X7 FLASH_ADC_SYM_4_0/a_200_531# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 FLASH_ADC_SYM_2_0/a_200_531# VIN GND GND sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X9 GND VIN FLASH_ADC_SYM_2_0/a_200_531# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X10 FLASH_ADC_SYM_2_0/a_200_531# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=3.528e+11p pd=3.08e+06u as=0p ps=0u w=1.26e+06u l=150000u
X11 T_2 FLASH_ADC_SYM_2_0/a_200_531# VDD VDD sky130_fd_pr__pfet_01v8 ad=3.528e+11p pd=3.08e+06u as=0p ps=0u w=1.26e+06u l=150000u
X12 VDD VIN FLASH_ADC_SYM_2_0/a_200_531# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X13 VDD FLASH_ADC_SYM_2_0/a_200_531# T_2 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.26e+06u l=150000u
X14 T_2 FLASH_ADC_SYM_2_0/a_200_531# GND GND sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X15 GND FLASH_ADC_SYM_2_0/a_200_531# T_2 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X16 FLASH_ADC_SYM_7_0/a_200_531# VIN GND GND sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X17 FLASH_ADC_SYM_7_0/a_200_531# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X18 T_7 FLASH_ADC_SYM_7_0/a_200_531# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X19 GND VIN FLASH_ADC_SYM_7_0/a_200_531# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X20 VDD VIN FLASH_ADC_SYM_7_0/a_200_531# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X21 VDD FLASH_ADC_SYM_7_0/a_200_531# T_7 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X22 T_7 FLASH_ADC_SYM_7_0/a_200_531# GND GND sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X23 GND FLASH_ADC_SYM_7_0/a_200_531# T_7 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X24 GND VIN FLASH_ADC_SYM_5_0/a_200_531# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.056e+11p ps=5.6e+06u w=2.52e+06u l=150000u
X25 FLASH_ADC_SYM_5_0/a_200_531# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X26 T_5 FLASH_ADC_SYM_5_0/a_200_531# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X27 VDD VIN FLASH_ADC_SYM_5_0/a_200_531# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X28 VDD FLASH_ADC_SYM_5_0/a_200_531# T_5 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X29 T_5 FLASH_ADC_SYM_5_0/a_200_531# GND GND sky130_fd_pr__nfet_01v8 ad=7.056e+11p pd=5.6e+06u as=0p ps=0u w=2.52e+06u l=150000u
X30 GND FLASH_ADC_SYM_5_0/a_200_531# T_5 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.52e+06u l=150000u
X31 FLASH_ADC_SYM_5_0/a_200_531# VIN GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.52e+06u l=150000u
X32 T_3 FLASH_ADC_SYM_3_0/a_200_531# GND GND sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X33 FLASH_ADC_SYM_3_0/a_200_531# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=0p ps=0u w=1.68e+06u l=150000u
X34 GND FLASH_ADC_SYM_3_0/a_200_531# T_3 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X35 T_3 FLASH_ADC_SYM_3_0/a_200_531# VDD VDD sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=0p ps=0u w=1.68e+06u l=150000u
X36 VDD VIN FLASH_ADC_SYM_3_0/a_200_531# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X37 VDD FLASH_ADC_SYM_3_0/a_200_531# T_3 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X38 FLASH_ADC_SYM_3_0/a_200_531# VIN GND GND sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X39 GND VIN FLASH_ADC_SYM_3_0/a_200_531# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X40 FLASH_ADC_SYM_1_0/a_200_531# VIN GND GND sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X41 GND VIN FLASH_ADC_SYM_1_0/a_200_531# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X42 FLASH_ADC_SYM_1_0/a_200_531# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=7.056e+11p pd=5.6e+06u as=0p ps=0u w=2.52e+06u l=150000u
X43 T_1 FLASH_ADC_SYM_1_0/a_200_531# VDD VDD sky130_fd_pr__pfet_01v8 ad=7.056e+11p pd=5.6e+06u as=0p ps=0u w=2.52e+06u l=150000u
X44 VDD VIN FLASH_ADC_SYM_1_0/a_200_531# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.52e+06u l=150000u
X45 VDD FLASH_ADC_SYM_1_0/a_200_531# T_1 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.52e+06u l=150000u
X46 T_1 FLASH_ADC_SYM_1_0/a_200_531# GND GND sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X47 GND FLASH_ADC_SYM_1_0/a_200_531# T_1 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X48 GND FLASH_ADC_SYM_6_0/a_200_531# T_6 GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.764e+11p ps=1.82e+06u w=630000u l=150000u
X49 FLASH_ADC_SYM_6_0/a_200_531# VIN VDD VDD sky130_fd_pr__pfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X50 T_6 FLASH_ADC_SYM_6_0/a_200_531# VDD VDD sky130_fd_pr__pfet_01v8 ad=1.176e+11p pd=1.4e+06u as=0p ps=0u w=420000u l=150000u
X51 VDD VIN FLASH_ADC_SYM_6_0/a_200_531# VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X52 FLASH_ADC_SYM_6_0/a_200_531# VIN GND GND sky130_fd_pr__nfet_01v8 ad=1.764e+11p pd=1.82e+06u as=0p ps=0u w=630000u l=150000u
X53 VDD FLASH_ADC_SYM_6_0/a_200_531# T_6 VDD sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
X54 GND VIN FLASH_ADC_SYM_6_0/a_200_531# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
X55 T_6 FLASH_ADC_SYM_6_0/a_200_531# GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=630000u l=150000u
C0 T_1 FLASH_ADC_SYM_7_0/a_200_531# 0.05fF
C1 FLASH_ADC_SYM_4_0/a_200_531# sky130_fd_sc_hd__fill_8_8/VPB 0.00fF
C2 VDD Y1 2.10fF
C3 sky130_fd_sc_hd__fill_2_7/VPB T_2 0.09fF
C4 T_6 T_2 0.33fF
C5 VDD sky130_fd_sc_hd__or4_1_0/a_277_297# 0.00fF
C6 Y2 sky130_fd_sc_hd__or4_1_1/a_27_297# 0.00fF
C7 T_3 T_5 0.21fF
C8 Y2 sky130_fd_sc_hd__or4_1_2/a_27_297# 0.02fF
C9 sky130_fd_sc_hd__fill_8_92/VPB GND 1.18fF
C10 T_6 sky130_fd_sc_hd__or4_1_1/a_277_297# 0.00fF
C11 T_3 T_7 0.44fF
C12 VDD sky130_fd_sc_hd__fill_8_8/VPB 1.64fF
C13 T_5 T_2 0.15fF
C14 sky130_fd_sc_hd__fill_8_93/VPB VDD 1.39fF
C15 T_7 T_2 0.12fF
C16 FLASH_ADC_SYM_6_0/a_200_531# VDD 2.93fF
C17 T_5 sky130_fd_sc_hd__or4_1_1/a_277_297# 0.00fF
C18 VDD FLASH_ADC_SYM_5_0/a_200_531# 3.17fF
C19 T_3 sky130_fd_sc_hd__or4_1_0/a_205_297# 0.00fF
C20 T_7 sky130_fd_sc_hd__or4_1_1/a_277_297# 0.00fF
C21 VIN T_3 0.51fF
C22 T_4 sky130_fd_sc_hd__or4_1_2/a_109_297# 0.00fF
C23 GND Y3 0.50fF
C24 Y2 sky130_fd_sc_hd__or4_1_2/a_277_297# 0.00fF
C25 Y2 sky130_fd_sc_hd__or4_1_0/a_27_297# 0.09fF
C26 Y1 sky130_fd_sc_hd__fill_2_7/VPB 0.03fF
C27 Y1 T_6 0.01fF
C28 VIN T_2 0.45fF
C29 T_4 T_1 0.08fF
C30 sky130_fd_sc_hd__or4_1_0/a_277_297# T_6 0.00fF
C31 Y1 T_5 0.12fF
C32 VDD Y2 3.12fF
C33 Y1 T_7 0.01fF
C34 sky130_fd_sc_hd__fill_8_93/VPB T_6 0.00fF
C35 sky130_fd_sc_hd__or4_1_0/a_277_297# T_7 0.00fF
C36 FLASH_ADC_SYM_6_0/a_200_531# T_6 0.39fF
C37 sky130_fd_sc_hd__fill_8_1/VPB T_3 0.00fF
C38 T_3 sky130_fd_sc_hd__fill_8_4/VPB 0.01fF
C39 T_6 FLASH_ADC_SYM_5_0/a_200_531# 0.30fF
C40 GND T_3 4.20fF
C41 sky130_fd_sc_hd__fill_8_1/VPB T_2 0.08fF
C42 T_2 sky130_fd_sc_hd__fill_8_4/VPB 0.07fF
C43 GND T_2 2.40fF
C44 FLASH_ADC_SYM_6_0/a_200_531# T_5 0.11fF
C45 T_5 FLASH_ADC_SYM_5_0/a_200_531# 0.47fF
C46 VIN Y1 0.07fF
C47 FLASH_ADC_SYM_6_0/a_200_531# T_7 0.00fF
C48 T_4 sky130_fd_sc_hd__or4_1_2/a_205_297# 0.00fF
C49 GND sky130_fd_sc_hd__or4_1_1/a_277_297# 0.00fF
C50 VIN sky130_fd_sc_hd__fill_8_8/VPB 0.34fF
C51 VDD FLASH_ADC_SYM_7_0/a_200_531# 2.95fF
C52 sky130_fd_sc_hd__or4_1_2/a_109_297# sky130_fd_sc_hd__or4_1_2/a_27_297# 0.02fF
C53 T_6 Y2 0.26fF
C54 sky130_fd_sc_hd__fill_8_87/VPB FLASH_ADC_SYM_5_0/a_200_531# 0.01fF
C55 T_4 sky130_fd_sc_hd__or4_1_2/a_27_297# 0.32fF
C56 FLASH_ADC_SYM_6_0/a_200_531# VIN 1.11fF
C57 T_1 sky130_fd_sc_hd__or4_1_1/a_27_297# 0.06fF
C58 VIN FLASH_ADC_SYM_5_0/a_200_531# 0.57fF
C59 T_5 Y2 0.00fF
C60 sky130_fd_sc_hd__fill_8_1/VPB Y1 0.02fF
C61 Y1 sky130_fd_sc_hd__fill_8_4/VPB 0.01fF
C62 GND Y1 2.13fF
C63 Y2 T_7 0.32fF
C64 GND sky130_fd_sc_hd__or4_1_0/a_277_297# 0.00fF
C65 GND sky130_fd_sc_hd__fill_8_8/VPB 1.40fF
C66 T_4 sky130_fd_sc_hd__or4_1_2/a_277_297# 0.00fF
C67 T_4 sky130_fd_sc_hd__or4_1_0/a_27_297# 0.00fF
C68 FLASH_ADC_SYM_4_0/a_200_531# T_4 0.26fF
C69 sky130_fd_sc_hd__fill_8_93/VPB GND 1.18fF
C70 FLASH_ADC_SYM_6_0/a_200_531# GND 0.06fF
C71 T_6 FLASH_ADC_SYM_7_0/a_200_531# 0.05fF
C72 sky130_fd_sc_hd__or4_1_2/a_205_297# sky130_fd_sc_hd__or4_1_2/a_27_297# 0.01fF
C73 VDD T_4 7.07fF
C74 T_5 FLASH_ADC_SYM_7_0/a_200_531# 0.11fF
C75 VDD T_1 5.19fF
C76 T_4 FLASH_ADC_SYM_3_0/a_200_531# 0.20fF
C77 T_3 T_2 3.00fF
C78 FLASH_ADC_SYM_7_0/a_200_531# T_7 0.37fF
C79 T_4 FLASH_ADC_SYM_2_0/a_200_531# 0.00fF
C80 sky130_fd_sc_hd__fill_8_92/VPB FLASH_ADC_SYM_5_0/a_200_531# 0.01fF
C81 T_3 sky130_fd_sc_hd__or4_1_1/a_277_297# 0.00fF
C82 GND Y2 0.56fF
C83 T_2 sky130_fd_sc_hd__or4_1_1/a_277_297# 0.00fF
C84 VIN FLASH_ADC_SYM_7_0/a_200_531# 0.96fF
C85 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_1/a_27_297# 0.01fF
C86 T_6 sky130_fd_sc_hd__or4_1_2/a_109_297# 0.00fF
C87 T_4 T_6 0.36fF
C88 sky130_fd_sc_hd__or4_1_2/a_277_297# sky130_fd_sc_hd__or4_1_2/a_27_297# 0.02fF
C89 FLASH_ADC_SYM_1_0/a_200_531# T_1 0.32fF
C90 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_2/a_27_297# 0.00fF
C91 T_3 Y1 1.41fF
C92 T_6 T_1 4.17fF
C93 T_5 sky130_fd_sc_hd__or4_1_2/a_109_297# 0.00fF
C94 T_4 T_5 0.47fF
C95 sky130_fd_sc_hd__or4_1_1/a_27_297# sky130_fd_sc_hd__or4_1_1/a_109_297# 0.02fF
C96 T_3 sky130_fd_sc_hd__or4_1_0/a_277_297# 0.00fF
C97 Y1 T_2 2.56fF
C98 T_7 sky130_fd_sc_hd__or4_1_2/a_109_297# 0.01fF
C99 VDD sky130_fd_sc_hd__or4_1_1/a_27_297# 0.27fF
C100 T_4 T_7 0.39fF
C101 sky130_fd_sc_hd__or4_1_0/a_277_297# T_2 0.00fF
C102 VDD sky130_fd_sc_hd__or4_1_2/a_27_297# 0.25fF
C103 T_5 T_1 1.30fF
C104 T_3 sky130_fd_sc_hd__fill_8_8/VPB 0.01fF
C105 Y1 sky130_fd_sc_hd__or4_1_1/a_277_297# 0.00fF
C106 GND FLASH_ADC_SYM_7_0/a_200_531# 0.02fF
C107 T_1 T_7 0.30fF
C108 sky130_fd_sc_hd__fill_8_8/VPB T_2 0.07fF
C109 Y2 Y3 1.66fF
C110 VIN T_4 1.00fF
C111 sky130_fd_sc_hd__fill_8_87/VPB T_1 0.11fF
C112 T_6 sky130_fd_sc_hd__or4_1_2/a_205_297# 0.00fF
C113 VDD sky130_fd_sc_hd__or4_1_2/a_277_297# 0.00fF
C114 VIN T_1 0.38fF
C115 VDD sky130_fd_sc_hd__or4_1_0/a_27_297# 0.36fF
C116 VDD FLASH_ADC_SYM_4_0/a_200_531# 2.90fF
C117 T_5 sky130_fd_sc_hd__or4_1_2/a_205_297# 0.00fF
C118 sky130_fd_sc_hd__or4_1_1/a_27_297# sky130_fd_sc_hd__or4_1_1/a_205_297# 0.01fF
C119 T_6 sky130_fd_sc_hd__or4_1_1/a_27_297# 0.03fF
C120 FLASH_ADC_SYM_4_0/a_200_531# FLASH_ADC_SYM_3_0/a_200_531# 0.00fF
C121 T_7 sky130_fd_sc_hd__or4_1_2/a_205_297# 0.00fF
C122 VDD sky130_fd_sc_hd__or4_1_1/a_109_297# 0.00fF
C123 T_6 sky130_fd_sc_hd__or4_1_2/a_27_297# 0.26fF
C124 T_3 Y2 0.11fF
C125 Y1 sky130_fd_sc_hd__fill_8_8/VPB 0.01fF
C126 T_5 sky130_fd_sc_hd__or4_1_1/a_27_297# 0.32fF
C127 GND sky130_fd_sc_hd__or4_1_2/a_109_297# 0.00fF
C128 Y2 T_2 0.01fF
C129 GND T_4 1.26fF
C130 T_5 sky130_fd_sc_hd__or4_1_2/a_27_297# 0.08fF
C131 T_7 sky130_fd_sc_hd__or4_1_1/a_27_297# 0.21fF
C132 VDD FLASH_ADC_SYM_3_0/a_200_531# 2.72fF
C133 T_7 sky130_fd_sc_hd__or4_1_2/a_27_297# 0.47fF
C134 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_0/a_109_297# 0.02fF
C135 GND T_1 2.99fF
C136 VDD FLASH_ADC_SYM_2_0/a_200_531# 2.87fF
C137 FLASH_ADC_SYM_3_0/a_200_531# FLASH_ADC_SYM_2_0/a_200_531# 0.00fF
C138 T_6 sky130_fd_sc_hd__or4_1_2/a_277_297# 0.00fF
C139 T_6 sky130_fd_sc_hd__or4_1_0/a_27_297# 0.22fF
C140 VDD sky130_fd_sc_hd__or4_1_0/a_109_297# 0.01fF
C141 sky130_fd_sc_hd__fill_8_93/VPB FLASH_ADC_SYM_5_0/a_200_531# 0.00fF
C142 T_5 sky130_fd_sc_hd__or4_1_2/a_277_297# 0.00fF
C143 VDD FLASH_ADC_SYM_1_0/a_200_531# 3.11fF
C144 FLASH_ADC_SYM_6_0/a_200_531# FLASH_ADC_SYM_5_0/a_200_531# 0.00fF
C145 T_5 sky130_fd_sc_hd__or4_1_0/a_27_297# 0.01fF
C146 T_6 sky130_fd_sc_hd__or4_1_1/a_109_297# 0.00fF
C147 FLASH_ADC_SYM_4_0/a_200_531# T_5 0.01fF
C148 sky130_fd_sc_hd__fill_8_92/VPB T_1 0.14fF
C149 T_7 sky130_fd_sc_hd__or4_1_2/a_277_297# 0.00fF
C150 VDD sky130_fd_sc_hd__or4_1_1/a_205_297# 0.00fF
C151 VDD sky130_fd_sc_hd__fill_2_7/VPB 1.31fF
C152 sky130_fd_sc_hd__or4_1_0/a_27_297# T_7 0.22fF
C153 VDD T_6 4.93fF
C154 T_5 sky130_fd_sc_hd__or4_1_1/a_109_297# 0.01fF
C155 sky130_fd_sc_hd__or4_1_0/a_277_297# Y2 0.00fF
C156 FLASH_ADC_SYM_1_0/a_200_531# FLASH_ADC_SYM_2_0/a_200_531# 0.00fF
C157 GND sky130_fd_sc_hd__or4_1_2/a_205_297# 0.00fF
C158 VDD T_5 5.05fF
C159 T_7 sky130_fd_sc_hd__or4_1_1/a_109_297# 0.00fF
C160 sky130_fd_sc_hd__or4_1_0/a_27_297# sky130_fd_sc_hd__or4_1_0/a_205_297# 0.01fF
C161 T_4 Y3 0.15fF
C162 VDD T_7 7.85fF
C163 T_5 FLASH_ADC_SYM_3_0/a_200_531# 0.02fF
C164 GND sky130_fd_sc_hd__or4_1_1/a_27_297# 0.36fF
C165 VIN FLASH_ADC_SYM_4_0/a_200_531# 1.11fF
C166 GND sky130_fd_sc_hd__or4_1_2/a_27_297# 0.36fF
C167 T_6 sky130_fd_sc_hd__or4_1_0/a_109_297# 0.00fF
C168 VDD sky130_fd_sc_hd__or4_1_0/a_205_297# 0.00fF
C169 VDD sky130_fd_sc_hd__fill_8_87/VPB 1.82fF
C170 VDD VIN 19.19fF
C171 T_5 sky130_fd_sc_hd__or4_1_0/a_109_297# 0.00fF
C172 T_6 sky130_fd_sc_hd__or4_1_1/a_205_297# 0.00fF
C173 sky130_fd_sc_hd__or4_1_0/a_109_297# T_7 0.00fF
C174 T_3 T_4 0.11fF
C175 VIN FLASH_ADC_SYM_3_0/a_200_531# 1.09fF
C176 T_2 sky130_fd_sc_hd__or4_1_2/a_109_297# 0.00fF
C177 T_5 sky130_fd_sc_hd__or4_1_1/a_205_297# 0.00fF
C178 T_4 T_2 0.08fF
C179 VIN FLASH_ADC_SYM_2_0/a_200_531# 1.18fF
C180 GND sky130_fd_sc_hd__or4_1_2/a_277_297# 0.00fF
C181 T_5 T_6 1.33fF
C182 T_3 T_1 0.00fF
C183 GND sky130_fd_sc_hd__or4_1_0/a_27_297# 0.28fF
C184 GND FLASH_ADC_SYM_4_0/a_200_531# 0.05fF
C185 T_7 sky130_fd_sc_hd__or4_1_1/a_205_297# 0.00fF
C186 T_6 T_7 0.87fF
C187 T_1 T_2 0.00fF
C188 FLASH_ADC_SYM_6_0/a_200_531# FLASH_ADC_SYM_7_0/a_200_531# 0.00fF
C189 GND sky130_fd_sc_hd__or4_1_1/a_109_297# 0.00fF
C190 T_5 T_7 1.77fF
C191 sky130_fd_sc_hd__fill_8_1/VPB VDD 1.89fF
C192 VDD sky130_fd_sc_hd__fill_8_4/VPB 1.25fF
C193 VDD GND 146.38fF
C194 T_6 sky130_fd_sc_hd__or4_1_0/a_205_297# 0.00fF
C195 FLASH_ADC_SYM_1_0/a_200_531# VIN 0.56fF
C196 sky130_fd_sc_hd__fill_8_87/VPB T_6 0.20fF
C197 Y3 sky130_fd_sc_hd__or4_1_2/a_27_297# 0.09fF
C198 VIN sky130_fd_sc_hd__fill_2_7/VPB 0.17fF
C199 GND FLASH_ADC_SYM_3_0/a_200_531# 0.06fF
C200 VIN T_6 0.42fF
C201 GND FLASH_ADC_SYM_2_0/a_200_531# 0.04fF
C202 T_5 sky130_fd_sc_hd__or4_1_0/a_205_297# 0.00fF
C203 Y1 T_4 0.00fF
C204 sky130_fd_sc_hd__or4_1_0/a_205_297# T_7 0.00fF
C205 VIN T_5 0.70fF
C206 sky130_fd_sc_hd__fill_8_92/VPB VDD 1.36fF
C207 VIN T_7 0.10fF
C208 Y1 T_1 0.00fF
C209 GND sky130_fd_sc_hd__or4_1_0/a_109_297# 0.00fF
C210 T_3 sky130_fd_sc_hd__or4_1_1/a_27_297# 0.23fF
C211 T_4 sky130_fd_sc_hd__fill_8_8/VPB 0.00fF
C212 Y3 sky130_fd_sc_hd__or4_1_2/a_277_297# 0.00fF
C213 FLASH_ADC_SYM_1_0/a_200_531# GND 0.15fF
C214 T_3 sky130_fd_sc_hd__or4_1_2/a_27_297# 0.00fF
C215 T_2 sky130_fd_sc_hd__or4_1_1/a_27_297# 0.01fF
C216 GND sky130_fd_sc_hd__or4_1_1/a_205_297# 0.00fF
C217 GND sky130_fd_sc_hd__fill_2_7/VPB 1.39fF
C218 VIN sky130_fd_sc_hd__fill_8_87/VPB 0.00fF
C219 T_2 sky130_fd_sc_hd__or4_1_2/a_27_297# 0.00fF
C220 GND T_6 5.50fF
C221 sky130_fd_sc_hd__fill_8_93/VPB T_1 0.11fF
C222 sky130_fd_sc_hd__or4_1_1/a_27_297# sky130_fd_sc_hd__or4_1_1/a_277_297# 0.01fF
C223 FLASH_ADC_SYM_6_0/a_200_531# T_1 0.05fF
C224 VDD Y3 0.64fF
C225 GND T_5 1.72fF
C226 T_1 FLASH_ADC_SYM_5_0/a_200_531# 0.10fF
C227 GND T_7 5.04fF
C228 T_3 sky130_fd_sc_hd__or4_1_0/a_27_297# 0.28fF
C229 T_3 FLASH_ADC_SYM_4_0/a_200_531# 0.09fF
C230 sky130_fd_sc_hd__fill_8_92/VPB T_6 0.05fF
C231 sky130_fd_sc_hd__or4_1_0/a_27_297# T_2 0.23fF
C232 FLASH_ADC_SYM_4_0/a_200_531# T_2 0.10fF
C233 GND sky130_fd_sc_hd__or4_1_0/a_205_297# 0.00fF
C234 GND sky130_fd_sc_hd__fill_8_87/VPB 1.17fF
C235 Y2 sky130_fd_sc_hd__or4_1_2/a_109_297# 0.00fF
C236 T_4 Y2 0.89fF
C237 T_3 sky130_fd_sc_hd__or4_1_1/a_109_297# 0.00fF
C238 Y1 sky130_fd_sc_hd__or4_1_1/a_27_297# 0.09fF
C239 sky130_fd_sc_hd__fill_8_92/VPB T_5 0.02fF
C240 sky130_fd_sc_hd__fill_8_1/VPB VIN 0.35fF
C241 VIN sky130_fd_sc_hd__fill_8_4/VPB 0.04fF
C242 VIN GND 6.71fF
C243 VDD T_3 4.60fF
C244 Y2 T_1 0.64fF
C245 VDD T_2 3.57fF
C246 T_3 FLASH_ADC_SYM_3_0/a_200_531# 0.34fF
C247 T_6 Y3 0.01fF
C248 T_3 FLASH_ADC_SYM_2_0/a_200_531# 0.24fF
C249 T_2 FLASH_ADC_SYM_3_0/a_200_531# 0.10fF
C250 VDD sky130_fd_sc_hd__or4_1_1/a_277_297# 0.00fF
C251 T_2 FLASH_ADC_SYM_2_0/a_200_531# 0.39fF
C252 T_5 Y3 0.00fF
C253 sky130_fd_sc_hd__fill_8_92/VPB VIN 0.00fF
C254 T_3 sky130_fd_sc_hd__or4_1_0/a_109_297# 0.00fF
C255 Y1 sky130_fd_sc_hd__or4_1_0/a_27_297# 0.00fF
C256 Y3 T_7 0.03fF
C257 sky130_fd_sc_hd__fill_8_1/VPB GND 1.25fF
C258 GND sky130_fd_sc_hd__fill_8_4/VPB 1.46fF
C259 Y1 FLASH_ADC_SYM_4_0/a_200_531# 0.00fF
C260 sky130_fd_sc_hd__or4_1_0/a_277_297# sky130_fd_sc_hd__or4_1_0/a_27_297# 0.01fF
C261 FLASH_ADC_SYM_1_0/a_200_531# T_3 0.00fF
C262 T_4 FLASH_ADC_SYM_7_0/a_200_531# 0.01fF
C263 Y2 sky130_fd_sc_hd__or4_1_2/a_205_297# 0.00fF
C264 T_3 sky130_fd_sc_hd__or4_1_1/a_205_297# 0.00fF
C265 T_3 sky130_fd_sc_hd__fill_2_7/VPB 0.00fF
C266 FLASH_ADC_SYM_1_0/a_200_531# T_2 0.00fF
C267 T_3 T_6 0.19fF
C268 VDD 0 217.43fF
C269 T_5 0 3.93fF
C270 Y1 0 3.10fF
C271 T_3 0 3.73fF
C272 GND 0 43.12fF
C273 T_2 0 3.03fF
C274 T_4 0 0.73fF
C275 Y3 0 2.17fF
C276 T_1 0 2.12fF
C277 Y2 0 0.55fF
C278 FLASH_ADC_SYM_6_0/a_200_531# 0 1.07fF
C279 sky130_fd_sc_hd__fill_8_93/VPB 0 4.35fF
C280 sky130_fd_sc_hd__fill_8_1/VPB 0 4.35fF
C281 sky130_fd_sc_hd__fill_8_8/VPB 0 4.35fF
C282 FLASH_ADC_SYM_1_0/a_200_531# 0 0.07fF
C283 FLASH_ADC_SYM_3_0/a_200_531# 0 0.59fF
C284 FLASH_ADC_SYM_5_0/a_200_531# 0 0.42fF
C285 FLASH_ADC_SYM_7_0/a_200_531# 0 1.10fF
C286 sky130_fd_sc_hd__fill_8_92/VPB 0 4.35fF
C287 sky130_fd_sc_hd__fill_8_4/VPB 0 4.35fF
C288 sky130_fd_sc_hd__fill_8_87/VPB 0 4.35fF
C289 sky130_fd_sc_hd__fill_2_7/VPB 0 4.35fF
C290 FLASH_ADC_SYM_2_0/a_200_531# 0 0.68fF
C291 FLASH_ADC_SYM_4_0/a_200_531# 0 0.53fF
.ends




*===============MANUALLY ADDED=========================
V1 VDD GND 1.8
.save i(v1)
V2 VIN GND sin(0 2 40Meg)
.save i(v2)
x1 T_1 T_6 T_7 VIN T_2 T_3 T_4 T_5 Y1 Y2 Y3 VDD GND flash_adc

**** begin user architecture code
.lib /home/swagatika/open_pdks/sky130/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.save all

.tran 0.001n 60n
.control
run
plot VIN VDD T_1 T_2 T_3 T_4 T_5 T_6 T_7
plot Y1 Y2+1.5 Y3+3
.save all
.endc
.end

**** end user architecture code
**.ends

