magic
tech sky130A
magscale 1 2
timestamp 1677569328
<< locali >>
rect 405 2419 413 2453
rect 447 2419 455 2453
rect 405 605 455 2419
rect 405 571 413 605
rect 447 571 455 605
<< viali >>
rect 413 2419 447 2453
rect 413 571 447 605
<< metal1 >>
rect 396 2453 464 2464
rect 396 2419 413 2453
rect 447 2419 464 2453
rect 396 2408 464 2419
rect 312 1622 376 1624
rect 312 1570 318 1622
rect 370 1570 376 1622
rect 312 1568 376 1570
rect 312 1454 376 1456
rect 312 1402 318 1454
rect 370 1402 376 1454
rect 312 1400 376 1402
rect 396 605 464 616
rect 396 571 413 605
rect 447 571 464 605
rect 396 560 464 571
<< via1 >>
rect 318 1570 370 1622
rect 318 1402 370 1454
<< metal2 >>
rect 316 1622 372 1628
rect 316 1570 318 1622
rect 370 1570 372 1622
rect 316 1454 372 1570
rect 316 1402 318 1454
rect 370 1402 372 1454
rect 316 1396 372 1402
use NMOS_S_21929916_X1_Y1_1677566905_1677566908  NMOS_S_21929916_X1_Y1_1677566905_1677566908_0
timestamp 1677569328
transform -1 0 516 0 -1 1512
box 52 56 395 1482
use PMOS_S_95864420_X1_Y1_1677566906_1677566908  PMOS_S_95864420_X1_Y1_1677566906_1677566908_0
timestamp 1677569328
transform -1 0 516 0 1 1512
box 0 0 516 1512
<< end >>
