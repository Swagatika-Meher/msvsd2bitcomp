VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Inverter_magic
  CLASS BLOCK ;
  FOREIGN Inverter_magic ;
  ORIGIN 6.000 6.370 ;
  SIZE 13.390 BY 15.550 ;
  PIN vdd
    ANTENNADIFFAREA 0.290000 ;
    PORT
      LAYER li1 ;
        RECT 0.485 3.810 0.655 4.850 ;
      LAYER mcon ;
        RECT 0.485 3.890 0.655 4.770 ;
      LAYER met1 ;
        RECT 0.280 7.760 1.280 9.180 ;
        RECT -2.460 6.930 1.280 7.760 ;
        RECT -2.440 6.460 1.280 6.930 ;
        RECT -2.440 4.820 -1.230 6.460 ;
        RECT 0.280 5.600 1.280 6.460 ;
        RECT 0.455 4.820 0.685 4.830 ;
        RECT -2.470 3.830 0.690 4.820 ;
    END
  END vdd
  PIN OUT
    ANTENNADIFFAREA 0.580000 ;
    PORT
      LAYER li1 ;
        RECT 0.925 3.810 1.095 4.850 ;
        RECT 0.920 -2.390 1.090 -1.350 ;
      LAYER mcon ;
        RECT 0.925 3.890 1.095 4.770 ;
        RECT 0.920 -2.310 1.090 -1.430 ;
      LAYER met1 ;
        RECT 0.920 4.830 3.580 4.840 ;
        RECT 0.895 3.830 4.440 4.830 ;
        RECT 0.920 3.800 4.440 3.830 ;
        RECT 3.120 1.360 4.440 3.800 ;
        RECT 3.120 0.370 7.390 1.360 ;
        RECT 3.120 -1.350 4.440 0.370 ;
        RECT 6.390 0.360 7.390 0.370 ;
        RECT 0.930 -1.370 4.440 -1.350 ;
        RECT 0.890 -2.370 4.440 -1.370 ;
        RECT 1.080 -2.390 4.440 -2.370 ;
    END
  END OUT
  PIN IN
    ANTENNAGATEAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT 0.625 5.065 0.955 5.235 ;
        RECT 0.625 3.425 0.955 3.595 ;
        RECT 0.620 -1.180 0.950 -1.010 ;
        RECT 0.620 -2.730 0.950 -2.560 ;
      LAYER mcon ;
        RECT 0.705 5.065 0.875 5.235 ;
        RECT 0.705 3.425 0.875 3.595 ;
        RECT 0.700 -1.180 0.870 -1.010 ;
        RECT 0.700 -2.730 0.870 -2.560 ;
      LAYER met1 ;
        RECT 0.630 5.030 0.940 5.290 ;
        RECT 0.630 5.020 0.930 5.030 ;
        RECT -1.910 3.660 0.780 3.680 ;
        RECT -1.910 3.650 0.860 3.660 ;
        RECT -2.460 3.625 0.860 3.650 ;
        RECT -2.460 3.395 0.935 3.625 ;
        RECT -2.460 3.340 0.860 3.395 ;
        RECT -6.000 1.340 -5.000 1.350 ;
        RECT -2.460 1.340 -1.340 3.340 ;
        RECT -6.000 0.350 -1.340 1.340 ;
        RECT -2.460 -0.920 -1.340 0.350 ;
        RECT -2.460 -0.980 0.920 -0.920 ;
        RECT -2.460 -1.210 0.930 -0.980 ;
        RECT -2.430 -1.220 0.790 -1.210 ;
        RECT 0.610 -2.800 0.940 -2.510 ;
    END
  END IN
  PIN gnd
    ANTENNADIFFAREA 0.290000 ;
    PORT
      LAYER li1 ;
        RECT 0.480 -2.390 0.650 -1.350 ;
      LAYER mcon ;
        RECT 0.480 -2.310 0.650 -1.430 ;
      LAYER met1 ;
        RECT 0.450 -1.410 0.680 -1.370 ;
        RECT -2.410 -1.430 0.680 -1.410 ;
        RECT -2.460 -2.360 0.680 -1.430 ;
        RECT -2.460 -3.940 -1.370 -2.360 ;
        RECT 0.450 -2.370 0.680 -2.360 ;
        RECT 0.280 -3.940 1.280 -3.060 ;
        RECT -2.460 -5.070 1.280 -3.940 ;
        RECT -2.440 -5.080 1.280 -5.070 ;
        RECT 0.280 -6.370 1.280 -5.080 ;
    END
  END gnd
  OBS
      LAYER nwell ;
        RECT -0.265 2.735 1.845 5.925 ;
      LAYER pwell ;
        RECT -0.270 -3.420 1.840 -0.320 ;
      LAYER li1 ;
        RECT -0.085 5.575 1.665 5.745 ;
        RECT -0.085 3.085 0.085 5.575 ;
        RECT 1.495 3.085 1.665 5.575 ;
        RECT -0.085 2.915 1.665 3.085 ;
        RECT -0.090 -0.670 1.660 -0.500 ;
        RECT -0.090 -3.070 0.080 -0.670 ;
        RECT 1.490 -3.070 1.660 -0.670 ;
        RECT -0.090 -3.240 1.660 -3.070 ;
  END
END Inverter_magic
END LIBRARY

