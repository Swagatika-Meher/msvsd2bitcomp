magic
tech sky130A
magscale 1 2
timestamp 1677569328
<< nwell >>
rect 0 0 688 1512
<< pmos >>
rect 200 462 230 672
rect 286 462 316 672
rect 372 462 402 672
rect 458 462 488 672
<< pdiff >>
rect 147 648 200 672
rect 147 614 155 648
rect 189 614 200 648
rect 147 580 200 614
rect 147 546 155 580
rect 189 546 200 580
rect 147 512 200 546
rect 147 478 155 512
rect 189 478 200 512
rect 147 462 200 478
rect 230 648 286 672
rect 230 614 241 648
rect 275 614 286 648
rect 230 580 286 614
rect 230 546 241 580
rect 275 546 286 580
rect 230 512 286 546
rect 230 478 241 512
rect 275 478 286 512
rect 230 462 286 478
rect 316 648 372 672
rect 316 614 327 648
rect 361 614 372 648
rect 316 580 372 614
rect 316 546 327 580
rect 361 546 372 580
rect 316 512 372 546
rect 316 478 327 512
rect 361 478 372 512
rect 316 462 372 478
rect 402 648 458 672
rect 402 614 413 648
rect 447 614 458 648
rect 402 580 458 614
rect 402 546 413 580
rect 447 546 458 580
rect 402 512 458 546
rect 402 478 413 512
rect 447 478 458 512
rect 402 462 458 478
rect 488 648 541 672
rect 488 614 499 648
rect 533 614 541 648
rect 488 580 541 614
rect 488 546 499 580
rect 533 546 541 580
rect 488 512 541 546
rect 488 478 499 512
rect 533 478 541 512
rect 488 462 541 478
<< pdiffc >>
rect 155 614 189 648
rect 155 546 189 580
rect 155 478 189 512
rect 241 614 275 648
rect 241 546 275 580
rect 241 478 275 512
rect 327 614 361 648
rect 327 546 361 580
rect 327 478 361 512
rect 413 614 447 648
rect 413 546 447 580
rect 413 478 447 512
rect 499 614 533 648
rect 499 546 533 580
rect 499 478 533 512
<< nsubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
rect 413 1361 447 1456
rect 413 1232 447 1327
<< nsubdiffcont >>
rect 241 1327 275 1361
rect 413 1327 447 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 672 230 897
rect 286 672 316 897
rect 372 941 488 951
rect 372 907 413 941
rect 447 907 488 941
rect 372 897 488 907
rect 372 672 402 897
rect 458 672 488 897
rect 200 252 230 462
rect 286 252 316 462
rect 372 252 402 462
rect 458 252 488 462
<< polycont >>
rect 241 907 275 941
rect 413 907 447 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 405 1361 455 1445
rect 405 1327 413 1361
rect 447 1327 455 1361
rect 405 1243 455 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 405 991 413 1025
rect 447 991 455 1025
rect 405 941 455 991
rect 405 907 413 941
rect 447 907 455 941
rect 405 823 455 907
rect 147 648 197 773
rect 147 614 155 648
rect 189 614 197 648
rect 147 580 197 614
rect 147 546 155 580
rect 189 546 197 580
rect 147 512 197 546
rect 147 478 155 512
rect 189 478 197 512
rect 147 269 197 478
rect 147 235 155 269
rect 189 235 197 269
rect 147 67 197 235
rect 233 648 283 773
rect 233 614 241 648
rect 275 614 283 648
rect 233 580 283 614
rect 233 546 241 580
rect 275 546 283 580
rect 233 512 283 546
rect 233 478 241 512
rect 275 478 283 512
rect 233 101 283 478
rect 233 67 241 101
rect 275 67 283 101
rect 319 648 369 773
rect 319 614 327 648
rect 361 614 369 648
rect 319 580 369 614
rect 319 546 327 580
rect 361 546 369 580
rect 319 512 369 546
rect 319 478 327 512
rect 361 478 369 512
rect 319 269 369 478
rect 319 235 327 269
rect 361 235 369 269
rect 319 67 369 235
rect 405 648 455 773
rect 405 614 413 648
rect 447 614 455 648
rect 405 580 455 614
rect 405 546 413 580
rect 447 546 455 580
rect 405 512 455 546
rect 405 478 413 512
rect 447 478 455 512
rect 405 185 455 478
rect 405 151 413 185
rect 447 151 455 185
rect 405 67 455 151
rect 491 648 541 773
rect 491 614 499 648
rect 533 614 541 648
rect 491 580 541 614
rect 491 546 499 580
rect 533 546 541 580
rect 491 512 541 546
rect 491 478 499 512
rect 533 478 541 512
rect 491 269 541 478
rect 491 235 499 269
rect 533 235 541 269
rect 491 67 541 235
<< viali >>
rect 241 1327 275 1361
rect 413 1327 447 1361
rect 241 907 275 941
rect 413 991 447 1025
rect 155 235 189 269
rect 241 67 275 101
rect 327 235 361 269
rect 413 151 447 185
rect 499 235 533 269
<< metal1 >>
rect 224 1370 550 1372
rect 224 1361 490 1370
rect 224 1327 241 1361
rect 275 1327 413 1361
rect 447 1327 490 1361
rect 224 1318 490 1327
rect 542 1318 550 1370
rect 224 1316 550 1318
rect 224 1025 464 1036
rect 224 991 413 1025
rect 447 991 464 1025
rect 224 980 464 991
rect 52 941 292 952
rect 52 907 241 941
rect 275 907 292 941
rect 52 896 292 907
rect 138 278 550 280
rect 138 269 490 278
rect 138 235 155 269
rect 189 235 327 269
rect 361 235 490 269
rect 138 226 490 235
rect 542 226 550 278
rect 138 224 550 226
rect 224 185 464 196
rect 224 151 413 185
rect 447 151 464 185
rect 224 140 464 151
rect 52 101 292 112
rect 52 67 241 101
rect 275 67 292 101
rect 52 56 292 67
<< via1 >>
rect 490 1318 542 1370
rect 490 269 542 278
rect 490 235 499 269
rect 499 235 533 269
rect 533 235 542 269
rect 490 226 542 235
<< metal2 >>
rect 488 1370 544 1376
rect 488 1318 490 1370
rect 542 1318 544 1370
rect 488 278 544 1318
rect 488 226 490 278
rect 542 226 544 278
rect 488 220 544 226
<< end >>
